magic
tech sky130A
magscale 1 2
timestamp 1655423120
<< metal1 >>
rect 235166 700408 235172 700460
rect 235224 700448 235230 700460
rect 305638 700448 305644 700460
rect 235224 700420 305644 700448
rect 235224 700408 235230 700420
rect 305638 700408 305644 700420
rect 305696 700408 305702 700460
rect 429838 700408 429844 700460
rect 429896 700448 429902 700460
rect 434714 700448 434720 700460
rect 429896 700420 434720 700448
rect 429896 700408 429902 700420
rect 434714 700408 434720 700420
rect 434772 700408 434778 700460
rect 170306 700340 170312 700392
rect 170364 700380 170370 700392
rect 434898 700380 434904 700392
rect 170364 700352 434904 700380
rect 170364 700340 170370 700352
rect 434898 700340 434904 700352
rect 434956 700340 434962 700392
rect 57790 700272 57796 700324
rect 57848 700312 57854 700324
rect 543458 700312 543464 700324
rect 57848 700284 543464 700312
rect 57848 700272 57854 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 147582 683136 147588 683188
rect 147640 683176 147646 683188
rect 580166 683176 580172 683188
rect 147640 683148 580172 683176
rect 147640 683136 147646 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 299474 640976 299480 641028
rect 299532 641016 299538 641028
rect 405734 641016 405740 641028
rect 299532 640988 405740 641016
rect 299532 640976 299538 640988
rect 405734 640976 405740 640988
rect 405792 640976 405798 641028
rect 104894 639548 104900 639600
rect 104952 639588 104958 639600
rect 434806 639588 434812 639600
rect 104952 639560 434812 639588
rect 104952 639548 104958 639560
rect 434806 639548 434812 639560
rect 434864 639548 434870 639600
rect 3418 638188 3424 638240
rect 3476 638228 3482 638240
rect 318150 638228 318156 638240
rect 3476 638200 318156 638228
rect 3476 638188 3482 638200
rect 318150 638188 318156 638200
rect 318208 638188 318214 638240
rect 364334 638188 364340 638240
rect 364392 638228 364398 638240
rect 428274 638228 428280 638240
rect 364392 638200 428280 638228
rect 364392 638188 364398 638200
rect 428274 638188 428280 638200
rect 428332 638188 428338 638240
rect 40034 636828 40040 636880
rect 40092 636868 40098 636880
rect 320818 636868 320824 636880
rect 40092 636840 320824 636868
rect 40092 636828 40098 636840
rect 320818 636828 320824 636840
rect 320876 636828 320882 636880
rect 307018 635740 307024 635792
rect 307076 635780 307082 635792
rect 355594 635780 355600 635792
rect 307076 635752 355600 635780
rect 307076 635740 307082 635752
rect 355594 635740 355600 635752
rect 355652 635740 355658 635792
rect 322474 635672 322480 635724
rect 322532 635712 322538 635724
rect 346578 635712 346584 635724
rect 322532 635684 346584 635712
rect 322532 635672 322538 635684
rect 346578 635672 346584 635684
rect 346636 635672 346642 635724
rect 322290 635604 322296 635656
rect 322348 635644 322354 635656
rect 432874 635644 432880 635656
rect 322348 635616 432880 635644
rect 322348 635604 322354 635616
rect 432874 635604 432880 635616
rect 432932 635604 432938 635656
rect 318058 635536 318064 635588
rect 318116 635576 318122 635588
rect 392302 635576 392308 635588
rect 318116 635548 392308 635576
rect 318116 635536 318122 635548
rect 392302 635536 392308 635548
rect 392360 635536 392366 635588
rect 323946 635468 323952 635520
rect 324004 635508 324010 635520
rect 369118 635508 369124 635520
rect 324004 635480 369124 635508
rect 324004 635468 324010 635480
rect 369118 635468 369124 635480
rect 369176 635468 369182 635520
rect 319438 635400 319444 635452
rect 319496 635440 319502 635452
rect 364610 635440 364616 635452
rect 319496 635412 364616 635440
rect 319496 635400 319502 635412
rect 364610 635400 364616 635412
rect 364668 635400 364674 635452
rect 316770 635332 316776 635384
rect 316828 635372 316834 635384
rect 342254 635372 342260 635384
rect 316828 635344 342260 635372
rect 316828 635332 316834 635344
rect 342254 635332 342260 635344
rect 342312 635332 342318 635384
rect 361390 635332 361396 635384
rect 361448 635372 361454 635384
rect 414842 635372 414848 635384
rect 361448 635344 414848 635372
rect 361448 635332 361454 635344
rect 414842 635332 414848 635344
rect 414900 635332 414906 635384
rect 324866 635264 324872 635316
rect 324924 635304 324930 635316
rect 378134 635304 378140 635316
rect 324924 635276 378140 635304
rect 324924 635264 324930 635276
rect 378134 635264 378140 635276
rect 378192 635264 378198 635316
rect 353294 635196 353300 635248
rect 353352 635236 353358 635248
rect 410334 635236 410340 635248
rect 353352 635208 410340 635236
rect 353352 635196 353358 635208
rect 410334 635196 410340 635208
rect 410392 635196 410398 635248
rect 313918 635128 313924 635180
rect 313976 635168 313982 635180
rect 373994 635168 374000 635180
rect 313976 635140 374000 635168
rect 313976 635128 313982 635140
rect 373994 635128 374000 635140
rect 374052 635128 374058 635180
rect 321002 635060 321008 635112
rect 321060 635100 321066 635112
rect 387794 635100 387800 635112
rect 321060 635072 387800 635100
rect 321060 635060 321066 635072
rect 387794 635060 387800 635072
rect 387852 635060 387858 635112
rect 314010 634992 314016 635044
rect 314068 635032 314074 635044
rect 383654 635032 383660 635044
rect 314068 635004 383660 635032
rect 314068 634992 314074 635004
rect 383654 634992 383660 635004
rect 383712 634992 383718 635044
rect 323854 634924 323860 634976
rect 323912 634964 323918 634976
rect 401594 634964 401600 634976
rect 323912 634936 401600 634964
rect 323912 634924 323918 634936
rect 401594 634924 401600 634936
rect 401652 634924 401658 634976
rect 322382 634856 322388 634908
rect 322440 634896 322446 634908
rect 337562 634896 337568 634908
rect 322440 634868 337568 634896
rect 322440 634856 322446 634868
rect 337562 634856 337568 634868
rect 337620 634856 337626 634908
rect 323762 634788 323768 634840
rect 323820 634828 323826 634840
rect 328638 634828 328644 634840
rect 323820 634800 328644 634828
rect 323820 634788 323826 634800
rect 328638 634788 328644 634800
rect 328696 634788 328702 634840
rect 391934 634788 391940 634840
rect 391992 634828 391998 634840
rect 419994 634828 420000 634840
rect 391992 634800 420000 634828
rect 391992 634788 391998 634800
rect 419994 634788 420000 634800
rect 420052 634828 420058 634840
rect 457438 634828 457444 634840
rect 420052 634800 457444 634828
rect 420052 634788 420058 634800
rect 457438 634788 457444 634800
rect 457496 634788 457502 634840
rect 323670 634312 323676 634364
rect 323728 634352 323734 634364
rect 436186 634352 436192 634364
rect 323728 634324 436192 634352
rect 323728 634312 323734 634324
rect 436186 634312 436192 634324
rect 436244 634312 436250 634364
rect 322566 634244 322572 634296
rect 322624 634284 322630 634296
rect 436094 634284 436100 634296
rect 322624 634256 436100 634284
rect 322624 634244 322630 634256
rect 436094 634244 436100 634256
rect 436152 634244 436158 634296
rect 236638 634176 236644 634228
rect 236696 634216 236702 634228
rect 360194 634216 360200 634228
rect 236696 634188 360200 634216
rect 236696 634176 236702 634188
rect 360194 634176 360200 634188
rect 360252 634176 360258 634228
rect 144914 634108 144920 634160
rect 144972 634148 144978 634160
rect 144972 634120 161474 634148
rect 144972 634108 144978 634120
rect 145006 634040 145012 634092
rect 145064 634080 145070 634092
rect 156598 634080 156604 634092
rect 145064 634052 156604 634080
rect 145064 634040 145070 634052
rect 156598 634040 156604 634052
rect 156656 634040 156662 634092
rect 161446 634080 161474 634120
rect 239398 634108 239404 634160
rect 239456 634148 239462 634160
rect 257062 634148 257068 634160
rect 239456 634120 257068 634148
rect 239456 634108 239462 634120
rect 257062 634108 257068 634120
rect 257120 634108 257126 634160
rect 322658 634108 322664 634160
rect 322716 634148 322722 634160
rect 457714 634148 457720 634160
rect 322716 634120 457720 634148
rect 322716 634108 322722 634120
rect 457714 634108 457720 634120
rect 457772 634108 457778 634160
rect 207658 634080 207664 634092
rect 161446 634052 207664 634080
rect 207658 634040 207664 634052
rect 207716 634040 207722 634092
rect 238202 634040 238208 634092
rect 238260 634080 238266 634092
rect 251358 634080 251364 634092
rect 238260 634052 251364 634080
rect 238260 634040 238266 634052
rect 251358 634040 251364 634052
rect 251416 634040 251422 634092
rect 324222 634040 324228 634092
rect 324280 634080 324286 634092
rect 494054 634080 494060 634092
rect 324280 634052 494060 634080
rect 324280 634040 324286 634052
rect 494054 634040 494060 634052
rect 494112 634040 494118 634092
rect 109954 633972 109960 634024
rect 110012 634012 110018 634024
rect 120902 634012 120908 634024
rect 110012 633984 120908 634012
rect 110012 633972 110018 633984
rect 120902 633972 120908 633984
rect 120960 633972 120966 634024
rect 148870 633972 148876 634024
rect 148928 634012 148934 634024
rect 172882 634012 172888 634024
rect 148928 633984 172888 634012
rect 148928 633972 148934 633984
rect 172882 633972 172888 633984
rect 172940 633972 172946 634024
rect 226334 633972 226340 634024
rect 226392 634012 226398 634024
rect 300302 634012 300308 634024
rect 226392 633984 300308 634012
rect 226392 633972 226398 633984
rect 300302 633972 300308 633984
rect 300360 633972 300366 634024
rect 316954 633972 316960 634024
rect 317012 634012 317018 634024
rect 457530 634012 457536 634024
rect 317012 633984 457536 634012
rect 317012 633972 317018 633984
rect 457530 633972 457536 633984
rect 457588 633972 457594 634024
rect 112530 633904 112536 633956
rect 112588 633944 112594 633956
rect 122926 633944 122932 633956
rect 112588 633916 122932 633944
rect 112588 633904 112594 633916
rect 122926 633904 122932 633916
rect 122984 633904 122990 633956
rect 140774 633904 140780 633956
rect 140832 633944 140838 633956
rect 167086 633944 167092 633956
rect 140832 633916 167092 633944
rect 140832 633904 140838 633916
rect 167086 633904 167092 633916
rect 167144 633904 167150 633956
rect 214006 633904 214012 633956
rect 214064 633944 214070 633956
rect 289262 633944 289268 633956
rect 214064 633916 289268 633944
rect 214064 633904 214070 633916
rect 289262 633904 289268 633916
rect 289320 633904 289326 633956
rect 314194 633904 314200 633956
rect 314252 633944 314258 633956
rect 456794 633944 456800 633956
rect 314252 633916 456800 633944
rect 314252 633904 314258 633916
rect 456794 633904 456800 633916
rect 456852 633904 456858 633956
rect 86770 633836 86776 633888
rect 86828 633876 86834 633888
rect 124306 633876 124312 633888
rect 86828 633848 124312 633876
rect 86828 633836 86834 633848
rect 124306 633836 124312 633848
rect 124364 633836 124370 633888
rect 148778 633836 148784 633888
rect 148836 633876 148842 633888
rect 176102 633876 176108 633888
rect 148836 633848 176108 633876
rect 148836 633836 148842 633848
rect 176102 633836 176108 633848
rect 176160 633836 176166 633888
rect 231118 633836 231124 633888
rect 231176 633876 231182 633888
rect 248782 633876 248788 633888
rect 231176 633848 248788 633876
rect 231176 633836 231182 633848
rect 248782 633836 248788 633848
rect 248840 633836 248846 633888
rect 304258 633836 304264 633888
rect 304316 633876 304322 633888
rect 457622 633876 457628 633888
rect 304316 633848 457628 633876
rect 304316 633836 304322 633848
rect 457622 633836 457628 633848
rect 457680 633836 457686 633888
rect 115658 633768 115664 633820
rect 115716 633808 115722 633820
rect 124582 633808 124588 633820
rect 115716 633780 124588 633808
rect 115716 633768 115722 633780
rect 124582 633768 124588 633780
rect 124640 633768 124646 633820
rect 149790 633768 149796 633820
rect 149848 633808 149854 633820
rect 190546 633808 190552 633820
rect 149848 633780 190552 633808
rect 149848 633768 149854 633780
rect 190546 633768 190552 633780
rect 190604 633768 190610 633820
rect 234614 633768 234620 633820
rect 234672 633808 234678 633820
rect 396810 633808 396816 633820
rect 234672 633780 396816 633808
rect 234672 633768 234678 633780
rect 396810 633768 396816 633780
rect 396868 633768 396874 633820
rect 106642 633700 106648 633752
rect 106700 633740 106706 633752
rect 120994 633740 121000 633752
rect 106700 633712 121000 633740
rect 106700 633700 106706 633712
rect 120994 633700 121000 633712
rect 121052 633700 121058 633752
rect 142154 633700 142160 633752
rect 142212 633740 142218 633752
rect 184474 633740 184480 633752
rect 142212 633712 184480 633740
rect 142212 633700 142218 633712
rect 184474 633700 184480 633712
rect 184532 633700 184538 633752
rect 239582 633700 239588 633752
rect 239640 633740 239646 633752
rect 274634 633740 274640 633752
rect 239640 633712 274640 633740
rect 239640 633700 239646 633712
rect 274634 633700 274640 633712
rect 274692 633700 274698 633752
rect 304350 633700 304356 633752
rect 304408 633740 304414 633752
rect 471606 633740 471612 633752
rect 304408 633712 471612 633740
rect 304408 633700 304414 633712
rect 471606 633700 471612 633712
rect 471664 633700 471670 633752
rect 56502 633632 56508 633684
rect 56560 633672 56566 633684
rect 77294 633672 77300 633684
rect 56560 633644 77300 633672
rect 56560 633632 56566 633644
rect 77294 633632 77300 633644
rect 77352 633632 77358 633684
rect 104066 633632 104072 633684
rect 104124 633672 104130 633684
rect 122190 633672 122196 633684
rect 104124 633644 122196 633672
rect 104124 633632 104130 633644
rect 122190 633632 122196 633644
rect 122248 633632 122254 633684
rect 156598 633632 156604 633684
rect 156656 633672 156662 633684
rect 196066 633672 196072 633684
rect 156656 633644 196072 633672
rect 156656 633632 156662 633644
rect 196066 633632 196072 633644
rect 196124 633632 196130 633684
rect 213914 633632 213920 633684
rect 213972 633672 213978 633684
rect 245654 633672 245660 633684
rect 213972 633644 245660 633672
rect 213972 633632 213978 633644
rect 245654 633632 245660 633644
rect 245712 633632 245718 633684
rect 249334 633632 249340 633684
rect 249392 633672 249398 633684
rect 295518 633672 295524 633684
rect 249392 633644 295524 633672
rect 249392 633632 249398 633644
rect 295518 633632 295524 633644
rect 295576 633632 295582 633684
rect 314102 633632 314108 633684
rect 314160 633672 314166 633684
rect 483198 633672 483204 633684
rect 314160 633644 483204 633672
rect 314160 633632 314166 633644
rect 483198 633632 483204 633644
rect 483256 633632 483262 633684
rect 55030 633564 55036 633616
rect 55088 633604 55094 633616
rect 80238 633604 80244 633616
rect 55088 633576 80244 633604
rect 55088 633564 55094 633576
rect 80238 633564 80244 633576
rect 80296 633564 80302 633616
rect 100662 633564 100668 633616
rect 100720 633604 100726 633616
rect 124490 633604 124496 633616
rect 100720 633576 124496 633604
rect 100720 633564 100726 633576
rect 124490 633564 124496 633576
rect 124548 633564 124554 633616
rect 147490 633564 147496 633616
rect 147548 633604 147554 633616
rect 199286 633604 199292 633616
rect 147548 633576 199292 633604
rect 147548 633564 147554 633576
rect 199286 633564 199292 633576
rect 199344 633564 199350 633616
rect 235258 633564 235264 633616
rect 235316 633604 235322 633616
rect 291838 633604 291844 633616
rect 235316 633576 291844 633604
rect 235316 633564 235322 633576
rect 291838 633564 291844 633576
rect 291896 633564 291902 633616
rect 322198 633564 322204 633616
rect 322256 633604 322262 633616
rect 494790 633604 494796 633616
rect 322256 633576 494796 633604
rect 322256 633564 322262 633576
rect 494790 633564 494796 633576
rect 494848 633564 494854 633616
rect 55122 633496 55128 633548
rect 55180 633536 55186 633548
rect 91830 633536 91836 633548
rect 55180 633508 91836 633536
rect 55180 633496 55186 633508
rect 91830 633496 91836 633508
rect 91888 633496 91894 633548
rect 95050 633496 95056 633548
rect 95108 633536 95114 633548
rect 121638 633536 121644 633548
rect 95108 633508 121644 633536
rect 95108 633496 95114 633508
rect 121638 633496 121644 633508
rect 121696 633496 121702 633548
rect 133874 633496 133880 633548
rect 133932 633536 133938 633548
rect 149974 633536 149980 633548
rect 133932 633508 149980 633536
rect 133932 633496 133938 633508
rect 149974 633496 149980 633508
rect 150032 633496 150038 633548
rect 201862 633536 201868 633548
rect 150084 633508 201868 633536
rect 54846 633428 54852 633480
rect 54904 633468 54910 633480
rect 88702 633468 88708 633480
rect 54904 633440 88708 633468
rect 54904 633428 54910 633440
rect 88702 633428 88708 633440
rect 88760 633428 88766 633480
rect 147398 633428 147404 633480
rect 147456 633468 147462 633480
rect 147456 633440 149652 633468
rect 147456 633428 147462 633440
rect 149624 633400 149652 633440
rect 149698 633428 149704 633480
rect 149756 633468 149762 633480
rect 150084 633468 150112 633508
rect 201862 633496 201868 633508
rect 201920 633496 201926 633548
rect 205542 633496 205548 633548
rect 205600 633536 205606 633548
rect 212626 633536 212632 633548
rect 205600 633508 212632 633536
rect 205600 633496 205606 633508
rect 212626 633496 212632 633508
rect 212684 633496 212690 633548
rect 237374 633496 237380 633548
rect 237432 633536 237438 633548
rect 254486 633536 254492 633548
rect 237432 633508 254492 633536
rect 237432 633496 237438 633508
rect 254486 633496 254492 633508
rect 254544 633496 254550 633548
rect 320910 633496 320916 633548
rect 320968 633536 320974 633548
rect 501230 633536 501236 633548
rect 320968 633508 501236 633536
rect 320968 633496 320974 633508
rect 501230 633496 501236 633508
rect 501288 633496 501294 633548
rect 164510 633468 164516 633480
rect 149756 633440 150112 633468
rect 150176 633440 164516 633468
rect 149756 633428 149762 633440
rect 150176 633400 150204 633440
rect 164510 633428 164516 633440
rect 164568 633428 164574 633480
rect 255314 633428 255320 633480
rect 255372 633468 255378 633480
rect 262950 633468 262956 633480
rect 255372 633440 262956 633468
rect 255372 633428 255378 633440
rect 262950 633428 262956 633440
rect 263008 633428 263014 633480
rect 316862 633428 316868 633480
rect 316920 633468 316926 633480
rect 512178 633468 512184 633480
rect 316920 633440 512184 633468
rect 316920 633428 316926 633440
rect 512178 633428 512184 633440
rect 512236 633428 512242 633480
rect 149624 633372 150204 633400
rect 223574 632952 223580 633004
rect 223632 632992 223638 633004
rect 249334 632992 249340 633004
rect 223632 632964 249340 632992
rect 223632 632952 223638 632964
rect 249334 632952 249340 632964
rect 249392 632952 249398 633004
rect 222194 632884 222200 632936
rect 222252 632924 222258 632936
rect 255314 632924 255320 632936
rect 222252 632896 255320 632924
rect 222252 632884 222258 632896
rect 255314 632884 255320 632896
rect 255372 632884 255378 632936
rect 3510 632816 3516 632868
rect 3568 632856 3574 632868
rect 353294 632856 353300 632868
rect 3568 632828 353300 632856
rect 3568 632816 3574 632828
rect 353294 632816 353300 632828
rect 353352 632816 353358 632868
rect 3602 632748 3608 632800
rect 3660 632788 3666 632800
rect 361390 632788 361396 632800
rect 3660 632760 361396 632788
rect 3660 632748 3666 632760
rect 361390 632748 361396 632760
rect 361448 632748 361454 632800
rect 237834 632680 237840 632732
rect 237892 632720 237898 632732
rect 391934 632720 391940 632732
rect 237892 632692 391940 632720
rect 237892 632680 237898 632692
rect 391934 632680 391940 632692
rect 391992 632680 391998 632732
rect 238938 632476 238944 632528
rect 238996 632516 239002 632528
rect 580166 632516 580172 632528
rect 238996 632488 580172 632516
rect 238996 632476 239002 632488
rect 580166 632476 580172 632488
rect 580224 632476 580230 632528
rect 3418 632408 3424 632460
rect 3476 632448 3482 632460
rect 323578 632448 323584 632460
rect 3476 632420 323584 632448
rect 3476 632408 3482 632420
rect 323578 632408 323584 632420
rect 323636 632408 323642 632460
rect 319622 632340 319628 632392
rect 319680 632380 319686 632392
rect 436278 632380 436284 632392
rect 319680 632352 436284 632380
rect 319680 632340 319686 632352
rect 436278 632340 436284 632352
rect 436336 632340 436342 632392
rect 239030 632272 239036 632324
rect 239088 632312 239094 632324
rect 433334 632312 433340 632324
rect 239088 632284 433340 632312
rect 239088 632272 239094 632284
rect 433334 632272 433340 632284
rect 433392 632272 433398 632324
rect 317046 632204 317052 632256
rect 317104 632244 317110 632256
rect 512086 632244 512092 632256
rect 317104 632216 512092 632244
rect 317104 632204 317110 632216
rect 512086 632204 512092 632216
rect 512144 632204 512150 632256
rect 319530 632136 319536 632188
rect 319588 632176 319594 632188
rect 511994 632176 512000 632188
rect 319588 632148 512000 632176
rect 319588 632136 319594 632148
rect 511994 632136 512000 632148
rect 512052 632136 512058 632188
rect 146110 631252 146116 631304
rect 146168 631292 146174 631304
rect 155494 631292 155500 631304
rect 146168 631264 155500 631292
rect 146168 631252 146174 631264
rect 155494 631252 155500 631264
rect 155552 631252 155558 631304
rect 228358 631252 228364 631304
rect 228416 631292 228422 631304
rect 280246 631292 280252 631304
rect 228416 631264 280252 631292
rect 228416 631252 228422 631264
rect 280246 631252 280252 631264
rect 280304 631252 280310 631304
rect 124858 631184 124864 631236
rect 124916 631224 124922 631236
rect 187694 631224 187700 631236
rect 124916 631196 187700 631224
rect 124916 631184 124922 631196
rect 187694 631184 187700 631196
rect 187752 631184 187758 631236
rect 233878 631184 233884 631236
rect 233936 631224 233942 631236
rect 266538 631224 266544 631236
rect 233936 631196 266544 631224
rect 233936 631184 233942 631196
rect 266538 631184 266544 631196
rect 266596 631184 266602 631236
rect 148962 631116 148968 631168
rect 149020 631156 149026 631168
rect 158714 631156 158720 631168
rect 149020 631128 158720 631156
rect 149020 631116 149026 631128
rect 158714 631116 158720 631128
rect 158772 631116 158778 631168
rect 238110 631116 238116 631168
rect 238168 631156 238174 631168
rect 277670 631156 277676 631168
rect 238168 631128 277676 631156
rect 238168 631116 238174 631128
rect 277670 631116 277676 631128
rect 277728 631116 277734 631168
rect 144178 631048 144184 631100
rect 144236 631088 144242 631100
rect 161474 631088 161480 631100
rect 144236 631060 161480 631088
rect 144236 631048 144242 631060
rect 161474 631048 161480 631060
rect 161532 631048 161538 631100
rect 231210 631048 231216 631100
rect 231268 631088 231274 631100
rect 271966 631088 271972 631100
rect 231268 631060 271972 631088
rect 231268 631048 231274 631060
rect 271966 631048 271972 631060
rect 272024 631048 272030 631100
rect 56410 630980 56416 631032
rect 56468 631020 56474 631032
rect 65518 631020 65524 631032
rect 56468 630992 65524 631020
rect 56468 630980 56474 630992
rect 65518 630980 65524 630992
rect 65576 630980 65582 631032
rect 149882 630980 149888 631032
rect 149940 631020 149946 631032
rect 170306 631020 170312 631032
rect 149940 630992 170312 631020
rect 149940 630980 149946 630992
rect 170306 630980 170312 630992
rect 170364 630980 170370 631032
rect 217318 630980 217324 631032
rect 217376 631020 217382 631032
rect 260374 631020 260380 631032
rect 217376 630992 260380 631020
rect 217376 630980 217382 630992
rect 260374 630980 260380 630992
rect 260432 630980 260438 631032
rect 56318 630912 56324 630964
rect 56376 630952 56382 630964
rect 71222 630952 71228 630964
rect 56376 630924 71228 630952
rect 56376 630912 56382 630924
rect 71222 630912 71228 630924
rect 71280 630912 71286 630964
rect 83458 630912 83464 630964
rect 83516 630952 83522 630964
rect 124398 630952 124404 630964
rect 83516 630924 124404 630952
rect 83516 630912 83522 630924
rect 124398 630912 124404 630924
rect 124456 630912 124462 630964
rect 136634 630912 136640 630964
rect 136692 630952 136698 630964
rect 178678 630952 178684 630964
rect 136692 630924 178684 630952
rect 136692 630912 136698 630924
rect 178678 630912 178684 630924
rect 178736 630912 178742 630964
rect 214558 630912 214564 630964
rect 214616 630952 214622 630964
rect 268654 630952 268660 630964
rect 214616 630924 268660 630952
rect 214616 630912 214622 630924
rect 268654 630912 268660 630924
rect 268712 630912 268718 630964
rect 59354 630844 59360 630896
rect 59412 630884 59418 630896
rect 97902 630884 97908 630896
rect 59412 630856 97908 630884
rect 59412 630844 59418 630856
rect 97902 630844 97908 630856
rect 97960 630844 97966 630896
rect 140038 630844 140044 630896
rect 140096 630884 140102 630896
rect 193490 630884 193496 630896
rect 140096 630856 193496 630884
rect 140096 630844 140102 630856
rect 193490 630844 193496 630856
rect 193548 630844 193554 630896
rect 220170 630844 220176 630896
rect 220228 630884 220234 630896
rect 283558 630884 283564 630896
rect 220228 630856 283564 630884
rect 220228 630844 220234 630856
rect 283558 630844 283564 630856
rect 283616 630844 283622 630896
rect 57698 630776 57704 630828
rect 57756 630816 57762 630828
rect 74626 630816 74632 630828
rect 57756 630788 74632 630816
rect 57756 630776 57762 630788
rect 74626 630776 74632 630788
rect 74684 630776 74690 630828
rect 124214 630776 124220 630828
rect 124272 630816 124278 630828
rect 182082 630816 182088 630828
rect 124272 630788 182088 630816
rect 124272 630776 124278 630788
rect 182082 630776 182088 630788
rect 182140 630776 182146 630828
rect 220078 630776 220084 630828
rect 220136 630816 220142 630828
rect 286134 630816 286140 630828
rect 220136 630788 286140 630816
rect 220136 630776 220142 630788
rect 286134 630776 286140 630788
rect 286192 630776 286198 630828
rect 54938 630708 54944 630760
rect 54996 630748 55002 630760
rect 62942 630748 62948 630760
rect 54996 630720 62948 630748
rect 54996 630708 55002 630720
rect 62942 630708 62948 630720
rect 63000 630708 63006 630760
rect 69290 630708 69296 630760
rect 69348 630748 69354 630760
rect 125778 630748 125784 630760
rect 69348 630720 125784 630748
rect 69348 630708 69354 630720
rect 125778 630708 125784 630720
rect 125836 630708 125842 630760
rect 148318 630708 148324 630760
rect 148376 630748 148382 630760
rect 153102 630748 153108 630760
rect 148376 630720 153108 630748
rect 148376 630708 148382 630720
rect 153102 630708 153108 630720
rect 153160 630708 153166 630760
rect 215938 630708 215944 630760
rect 215996 630748 216002 630760
rect 297726 630748 297732 630760
rect 215996 630720 297732 630748
rect 215996 630708 216002 630720
rect 297726 630708 297732 630720
rect 297784 630708 297790 630760
rect 57882 630640 57888 630692
rect 57940 630680 57946 630692
rect 146202 630680 146208 630692
rect 57940 630652 146208 630680
rect 57940 630640 57946 630652
rect 146202 630640 146208 630652
rect 146260 630680 146266 630692
rect 237834 630680 237840 630692
rect 146260 630652 237840 630680
rect 146260 630640 146266 630652
rect 237834 630640 237840 630652
rect 237892 630640 237898 630692
rect 239490 630640 239496 630692
rect 239548 630680 239554 630692
rect 242894 630680 242900 630692
rect 239548 630652 242900 630680
rect 239548 630640 239554 630652
rect 242894 630640 242900 630652
rect 242952 630640 242958 630692
rect 118142 630368 118148 630420
rect 118200 630408 118206 630420
rect 121454 630408 121460 630420
rect 118200 630380 121460 630408
rect 118200 630368 118206 630380
rect 121454 630368 121460 630380
rect 121512 630368 121518 630420
rect 215294 629892 215300 629944
rect 215352 629932 215358 629944
rect 237374 629932 237380 629944
rect 215352 629904 237380 629932
rect 215352 629892 215358 629904
rect 237374 629892 237380 629904
rect 237432 629892 237438 629944
rect 144270 627920 144276 627972
rect 144328 627960 144334 627972
rect 146294 627960 146300 627972
rect 144328 627932 146300 627960
rect 144328 627920 144334 627932
rect 146294 627920 146300 627932
rect 146352 627920 146358 627972
rect 217410 627920 217416 627972
rect 217468 627960 217474 627972
rect 237374 627960 237380 627972
rect 217468 627932 237380 627960
rect 217468 627920 217474 627932
rect 237374 627920 237380 627932
rect 237432 627920 237438 627972
rect 465442 627920 465448 627972
rect 465500 627960 465506 627972
rect 580258 627960 580264 627972
rect 465500 627932 580264 627960
rect 465500 627920 465506 627932
rect 580258 627920 580264 627932
rect 580316 627920 580322 627972
rect 238846 627784 238852 627836
rect 238904 627824 238910 627836
rect 239766 627824 239772 627836
rect 238904 627796 239772 627824
rect 238904 627784 238910 627796
rect 239766 627784 239772 627796
rect 239824 627784 239830 627836
rect 309778 626560 309784 626612
rect 309836 626600 309842 626612
rect 321554 626600 321560 626612
rect 309836 626572 321560 626600
rect 309836 626560 309842 626572
rect 321554 626560 321560 626572
rect 321612 626560 321618 626612
rect 233234 622412 233240 622464
rect 233292 622452 233298 622464
rect 237374 622452 237380 622464
rect 233292 622424 237380 622452
rect 233292 622412 233298 622424
rect 237374 622412 237380 622424
rect 237432 622412 237438 622464
rect 311158 622412 311164 622464
rect 311216 622452 311222 622464
rect 321554 622452 321560 622464
rect 311216 622424 321560 622452
rect 311216 622412 311222 622424
rect 321554 622412 321560 622424
rect 321612 622412 321618 622464
rect 140866 619624 140872 619676
rect 140924 619664 140930 619676
rect 146294 619664 146300 619676
rect 140924 619636 146300 619664
rect 140924 619624 140930 619636
rect 146294 619624 146300 619636
rect 146352 619624 146358 619676
rect 232498 619624 232504 619676
rect 232556 619664 232562 619676
rect 237374 619664 237380 619676
rect 232556 619636 237380 619664
rect 232556 619624 232562 619636
rect 237374 619624 237380 619636
rect 237432 619624 237438 619676
rect 316678 616836 316684 616888
rect 316736 616876 316742 616888
rect 321554 616876 321560 616888
rect 316736 616848 321560 616876
rect 316736 616836 316742 616848
rect 321554 616836 321560 616848
rect 321612 616836 321618 616888
rect 132494 615476 132500 615528
rect 132552 615516 132558 615528
rect 146294 615516 146300 615528
rect 132552 615488 146300 615516
rect 132552 615476 132558 615488
rect 146294 615476 146300 615488
rect 146352 615476 146358 615528
rect 222838 615476 222844 615528
rect 222896 615516 222902 615528
rect 237374 615516 237380 615528
rect 222896 615488 237380 615516
rect 222896 615476 222902 615488
rect 237374 615476 237380 615488
rect 237432 615476 237438 615528
rect 223666 612756 223672 612808
rect 223724 612796 223730 612808
rect 237374 612796 237380 612808
rect 223724 612768 237380 612796
rect 223724 612756 223730 612768
rect 237374 612756 237380 612768
rect 237432 612756 237438 612808
rect 312538 612756 312544 612808
rect 312596 612796 312602 612808
rect 321554 612796 321560 612808
rect 312596 612768 321560 612796
rect 312596 612756 312602 612768
rect 321554 612756 321560 612768
rect 321612 612756 321618 612808
rect 218054 609968 218060 610020
rect 218112 610008 218118 610020
rect 237374 610008 237380 610020
rect 218112 609980 237380 610008
rect 218112 609968 218118 609980
rect 237374 609968 237380 609980
rect 237432 609968 237438 610020
rect 312630 607180 312636 607232
rect 312688 607220 312694 607232
rect 321554 607220 321560 607232
rect 312688 607192 321560 607220
rect 312688 607180 312694 607192
rect 321554 607180 321560 607192
rect 321612 607180 321618 607232
rect 307110 603100 307116 603152
rect 307168 603140 307174 603152
rect 321554 603140 321560 603152
rect 307168 603112 321560 603140
rect 307168 603100 307174 603112
rect 321554 603100 321560 603112
rect 321612 603100 321618 603152
rect 229738 600312 229744 600364
rect 229796 600352 229802 600364
rect 237374 600352 237380 600364
rect 229796 600324 237380 600352
rect 229796 600312 229802 600324
rect 237374 600312 237380 600324
rect 237432 600312 237438 600364
rect 128998 597524 129004 597576
rect 129056 597564 129062 597576
rect 146294 597564 146300 597576
rect 129056 597536 146300 597564
rect 129056 597524 129062 597536
rect 146294 597524 146300 597536
rect 146352 597524 146358 597576
rect 217502 597524 217508 597576
rect 217560 597564 217566 597576
rect 237374 597564 237380 597576
rect 217560 597536 237380 597564
rect 217560 597524 217566 597536
rect 237374 597524 237380 597536
rect 237432 597524 237438 597576
rect 307202 597524 307208 597576
rect 307260 597564 307266 597576
rect 321554 597564 321560 597576
rect 307260 597536 321560 597564
rect 307260 597524 307266 597536
rect 321554 597524 321560 597536
rect 321612 597524 321618 597576
rect 302694 596776 302700 596828
rect 302752 596816 302758 596828
rect 322658 596816 322664 596828
rect 302752 596788 322664 596816
rect 302752 596776 302758 596788
rect 322658 596776 322664 596788
rect 322716 596776 322722 596828
rect 124122 596164 124128 596216
rect 124180 596204 124186 596216
rect 145558 596204 145564 596216
rect 124180 596176 145564 596204
rect 124180 596164 124186 596176
rect 145558 596164 145564 596176
rect 145616 596164 145622 596216
rect 214650 594804 214656 594856
rect 214708 594844 214714 594856
rect 237374 594844 237380 594856
rect 214708 594816 237380 594844
rect 214708 594804 214714 594816
rect 237374 594804 237380 594816
rect 237432 594804 237438 594856
rect 57422 591336 57428 591388
rect 57480 591376 57486 591388
rect 58618 591376 58624 591388
rect 57480 591348 58624 591376
rect 57480 591336 57486 591348
rect 58618 591336 58624 591348
rect 58676 591336 58682 591388
rect 220262 590656 220268 590708
rect 220320 590696 220326 590708
rect 237374 590696 237380 590708
rect 220320 590668 237380 590696
rect 220320 590656 220326 590668
rect 237374 590656 237380 590668
rect 237432 590656 237438 590708
rect 305730 589296 305736 589348
rect 305788 589336 305794 589348
rect 321554 589336 321560 589348
rect 305788 589308 321560 589336
rect 305788 589296 305794 589308
rect 321554 589296 321560 589308
rect 321612 589296 321618 589348
rect 231854 587868 231860 587920
rect 231912 587908 231918 587920
rect 237374 587908 237380 587920
rect 231912 587880 237380 587908
rect 231912 587868 231918 587880
rect 237374 587868 237380 587880
rect 237432 587868 237438 587920
rect 125594 585148 125600 585200
rect 125652 585188 125658 585200
rect 146294 585188 146300 585200
rect 125652 585160 146300 585188
rect 125652 585148 125658 585160
rect 146294 585148 146300 585160
rect 146352 585148 146358 585200
rect 235350 585148 235356 585200
rect 235408 585188 235414 585200
rect 237374 585188 237380 585200
rect 235408 585160 237380 585188
rect 235408 585148 235414 585160
rect 237374 585148 237380 585160
rect 237432 585148 237438 585200
rect 307294 583720 307300 583772
rect 307352 583760 307358 583772
rect 321554 583760 321560 583772
rect 307352 583732 321560 583760
rect 307352 583720 307358 583732
rect 321554 583720 321560 583732
rect 321612 583720 321618 583772
rect 130378 582360 130384 582412
rect 130436 582400 130442 582412
rect 146294 582400 146300 582412
rect 130436 582372 146300 582400
rect 130436 582360 130442 582372
rect 146294 582360 146300 582372
rect 146352 582360 146358 582412
rect 57790 581612 57796 581664
rect 57848 581652 57854 581664
rect 58710 581652 58716 581664
rect 57848 581624 58716 581652
rect 57848 581612 57854 581624
rect 58710 581612 58716 581624
rect 58768 581612 58774 581664
rect 139394 579640 139400 579692
rect 139452 579680 139458 579692
rect 146294 579680 146300 579692
rect 139452 579652 146300 579680
rect 139452 579640 139458 579652
rect 146294 579640 146300 579652
rect 146352 579640 146358 579692
rect 216030 579640 216036 579692
rect 216088 579680 216094 579692
rect 237374 579680 237380 579692
rect 216088 579652 237380 579680
rect 216088 579640 216094 579652
rect 237374 579640 237380 579652
rect 237432 579640 237438 579692
rect 317138 579640 317144 579692
rect 317196 579680 317202 579692
rect 321554 579680 321560 579692
rect 317196 579652 321560 579680
rect 317196 579640 317202 579652
rect 321554 579640 321560 579652
rect 321612 579640 321618 579692
rect 513006 579640 513012 579692
rect 513064 579680 513070 579692
rect 560938 579680 560944 579692
rect 513064 579652 560944 579680
rect 513064 579640 513070 579652
rect 560938 579640 560944 579652
rect 560996 579640 561002 579692
rect 226426 576852 226432 576904
rect 226484 576892 226490 576904
rect 237374 576892 237380 576904
rect 226484 576864 237380 576892
rect 226484 576852 226490 576864
rect 237374 576852 237380 576864
rect 237432 576852 237438 576904
rect 311250 574064 311256 574116
rect 311308 574104 311314 574116
rect 321554 574104 321560 574116
rect 311308 574076 321560 574104
rect 311308 574064 311314 574076
rect 321554 574064 321560 574076
rect 321612 574064 321618 574116
rect 218146 572704 218152 572756
rect 218204 572744 218210 572756
rect 237374 572744 237380 572756
rect 218204 572716 237380 572744
rect 218204 572704 218210 572716
rect 237374 572704 237380 572716
rect 237432 572704 237438 572756
rect 220354 569916 220360 569968
rect 220412 569956 220418 569968
rect 237374 569956 237380 569968
rect 220412 569928 237380 569956
rect 220412 569916 220418 569928
rect 237374 569916 237380 569928
rect 237432 569916 237438 569968
rect 318150 569848 318156 569900
rect 318208 569888 318214 569900
rect 321554 569888 321560 569900
rect 318208 569860 321560 569888
rect 318208 569848 318214 569860
rect 321554 569848 321560 569860
rect 321612 569848 321618 569900
rect 57146 569168 57152 569220
rect 57204 569208 57210 569220
rect 59906 569208 59912 569220
rect 57204 569180 59912 569208
rect 57204 569168 57210 569180
rect 59906 569168 59912 569180
rect 59964 569168 59970 569220
rect 3418 568488 3424 568540
rect 3476 568528 3482 568540
rect 307294 568528 307300 568540
rect 3476 568500 307300 568528
rect 3476 568488 3482 568500
rect 307294 568488 307300 568500
rect 307352 568488 307358 568540
rect 57330 568420 57336 568472
rect 57388 568460 57394 568472
rect 60734 568460 60740 568472
rect 57388 568432 60740 568460
rect 57388 568420 57394 568432
rect 60734 568420 60740 568432
rect 60792 568420 60798 568472
rect 113174 568420 113180 568472
rect 113232 568460 113238 568472
rect 122282 568460 122288 568472
rect 113232 568432 122288 568460
rect 113232 568420 113238 568432
rect 122282 568420 122288 568432
rect 122340 568420 122346 568472
rect 145558 568420 145564 568472
rect 145616 568460 145622 568472
rect 214098 568460 214104 568472
rect 145616 568432 214104 568460
rect 145616 568420 145622 568432
rect 214098 568420 214104 568432
rect 214156 568460 214162 568472
rect 302694 568460 302700 568472
rect 214156 568432 302700 568460
rect 214156 568420 214162 568432
rect 302694 568420 302700 568432
rect 302752 568420 302758 568472
rect 106274 568352 106280 568404
rect 106332 568392 106338 568404
rect 124582 568392 124588 568404
rect 106332 568364 124588 568392
rect 106332 568352 106338 568364
rect 124582 568352 124588 568364
rect 124640 568352 124646 568404
rect 147122 568352 147128 568404
rect 147180 568392 147186 568404
rect 151078 568392 151084 568404
rect 147180 568364 151084 568392
rect 147180 568352 147186 568364
rect 151078 568352 151084 568364
rect 151136 568352 151142 568404
rect 288526 568352 288532 568404
rect 288584 568392 288590 568404
rect 316862 568392 316868 568404
rect 288584 568364 316868 568392
rect 288584 568352 288590 568364
rect 316862 568352 316868 568364
rect 316920 568352 316926 568404
rect 99558 568284 99564 568336
rect 99616 568324 99622 568336
rect 123570 568324 123576 568336
rect 99616 568296 123576 568324
rect 99616 568284 99622 568296
rect 123570 568284 123576 568296
rect 123628 568284 123634 568336
rect 288618 568284 288624 568336
rect 288676 568324 288682 568336
rect 316954 568324 316960 568336
rect 288676 568296 316960 568324
rect 288676 568284 288682 568296
rect 316954 568284 316960 568296
rect 317012 568284 317018 568336
rect 96706 568216 96712 568268
rect 96764 568256 96770 568268
rect 122926 568256 122932 568268
rect 96764 568228 122932 568256
rect 96764 568216 96770 568228
rect 122926 568216 122932 568228
rect 122984 568216 122990 568268
rect 287054 568216 287060 568268
rect 287112 568256 287118 568268
rect 317046 568256 317052 568268
rect 287112 568228 317052 568256
rect 287112 568216 287118 568228
rect 317046 568216 317052 568228
rect 317104 568216 317110 568268
rect 87046 568148 87052 568200
rect 87104 568188 87110 568200
rect 121362 568188 121368 568200
rect 87104 568160 121368 568188
rect 87104 568148 87110 568160
rect 121362 568148 121368 568160
rect 121420 568148 121426 568200
rect 149698 568148 149704 568200
rect 149756 568188 149762 568200
rect 154758 568188 154764 568200
rect 149756 568160 154764 568188
rect 149756 568148 149762 568160
rect 154758 568148 154764 568160
rect 154816 568148 154822 568200
rect 204898 568148 204904 568200
rect 204956 568188 204962 568200
rect 212902 568188 212908 568200
rect 204956 568160 212908 568188
rect 204956 568148 204962 568160
rect 212902 568148 212908 568160
rect 212960 568148 212966 568200
rect 266354 568148 266360 568200
rect 266412 568188 266418 568200
rect 314010 568188 314016 568200
rect 266412 568160 314016 568188
rect 266412 568148 266418 568160
rect 314010 568148 314016 568160
rect 314068 568148 314074 568200
rect 58802 568080 58808 568132
rect 58860 568120 58866 568132
rect 67634 568120 67640 568132
rect 58860 568092 67640 568120
rect 58860 568080 58866 568092
rect 67634 568080 67640 568092
rect 67692 568080 67698 568132
rect 93854 568080 93860 568132
rect 93912 568120 93918 568132
rect 124490 568120 124496 568132
rect 93912 568092 124496 568120
rect 93912 568080 93918 568092
rect 124490 568080 124496 568092
rect 124548 568080 124554 568132
rect 147490 568080 147496 568132
rect 147548 568120 147554 568132
rect 156046 568120 156052 568132
rect 147548 568092 156052 568120
rect 147548 568080 147554 568092
rect 156046 568080 156052 568092
rect 156104 568080 156110 568132
rect 164418 568080 164424 568132
rect 164476 568120 164482 568132
rect 212626 568120 212632 568132
rect 164476 568092 212632 568120
rect 164476 568080 164482 568092
rect 212626 568080 212632 568092
rect 212684 568080 212690 568132
rect 260834 568080 260840 568132
rect 260892 568120 260898 568132
rect 319622 568120 319628 568132
rect 260892 568092 319628 568120
rect 260892 568080 260898 568092
rect 319622 568080 319628 568092
rect 319680 568080 319686 568132
rect 58986 568012 58992 568064
rect 59044 568052 59050 568064
rect 74534 568052 74540 568064
rect 59044 568024 74540 568052
rect 59044 568012 59050 568024
rect 74534 568012 74540 568024
rect 74592 568012 74598 568064
rect 98086 568012 98092 568064
rect 98144 568052 98150 568064
rect 120902 568052 120908 568064
rect 98144 568024 120908 568052
rect 98144 568012 98150 568024
rect 120902 568012 120908 568024
rect 120960 568012 120966 568064
rect 121454 568012 121460 568064
rect 121512 568052 121518 568064
rect 211246 568052 211252 568064
rect 121512 568024 211252 568052
rect 121512 568012 121518 568024
rect 211246 568012 211252 568024
rect 211304 568012 211310 568064
rect 258074 568012 258080 568064
rect 258132 568052 258138 568064
rect 322566 568052 322572 568064
rect 258132 568024 322572 568052
rect 258132 568012 258138 568024
rect 322566 568012 322572 568024
rect 322624 568012 322630 568064
rect 54846 567944 54852 567996
rect 54904 567984 54910 567996
rect 78674 567984 78680 567996
rect 54904 567956 78680 567984
rect 54904 567944 54910 567956
rect 78674 567944 78680 567956
rect 78732 567944 78738 567996
rect 86954 567944 86960 567996
rect 87012 567984 87018 567996
rect 120994 567984 121000 567996
rect 87012 567956 121000 567984
rect 87012 567944 87018 567956
rect 120994 567944 121000 567956
rect 121052 567944 121058 567996
rect 147398 567944 147404 567996
rect 147456 567984 147462 567996
rect 157334 567984 157340 567996
rect 147456 567956 157340 567984
rect 147456 567944 147462 567956
rect 157334 567944 157340 567956
rect 157392 567944 157398 567996
rect 194778 567944 194784 567996
rect 194836 567984 194842 567996
rect 302326 567984 302332 567996
rect 194836 567956 302332 567984
rect 194836 567944 194842 567956
rect 302326 567944 302332 567956
rect 302384 567944 302390 567996
rect 66346 567876 66352 567928
rect 66404 567916 66410 567928
rect 121546 567916 121552 567928
rect 66404 567888 121552 567916
rect 66404 567876 66410 567888
rect 121546 567876 121552 567888
rect 121604 567876 121610 567928
rect 148778 567876 148784 567928
rect 148836 567916 148842 567928
rect 161474 567916 161480 567928
rect 148836 567888 161480 567916
rect 148836 567876 148842 567888
rect 161474 567876 161480 567888
rect 161532 567876 161538 567928
rect 183646 567876 183652 567928
rect 183704 567916 183710 567928
rect 301130 567916 301136 567928
rect 183704 567888 301136 567916
rect 183704 567876 183710 567888
rect 301130 567876 301136 567888
rect 301188 567876 301194 567928
rect 63494 567808 63500 567860
rect 63552 567848 63558 567860
rect 123478 567848 123484 567860
rect 63552 567820 123484 567848
rect 63552 567808 63558 567820
rect 123478 567808 123484 567820
rect 123536 567808 123542 567860
rect 148870 567808 148876 567860
rect 148928 567848 148934 567860
rect 164326 567848 164332 567860
rect 148928 567820 164332 567848
rect 148928 567808 148934 567820
rect 164326 567808 164332 567820
rect 164384 567808 164390 567860
rect 179414 567808 179420 567860
rect 179472 567848 179478 567860
rect 300854 567848 300860 567860
rect 179472 567820 300860 567848
rect 179472 567808 179478 567820
rect 300854 567808 300860 567820
rect 300912 567808 300918 567860
rect 293954 567740 293960 567792
rect 294012 567780 294018 567792
rect 319530 567780 319536 567792
rect 294012 567752 319536 567780
rect 294012 567740 294018 567752
rect 319530 567740 319536 567752
rect 319588 567740 319594 567792
rect 289814 567672 289820 567724
rect 289872 567712 289878 567724
rect 314102 567712 314108 567724
rect 289872 567684 314108 567712
rect 289872 567672 289878 567684
rect 314102 567672 314108 567684
rect 314160 567672 314166 567724
rect 291194 567604 291200 567656
rect 291252 567644 291258 567656
rect 314194 567644 314200 567656
rect 291252 567616 314200 567644
rect 291252 567604 291258 567616
rect 314194 567604 314200 567616
rect 314252 567604 314258 567656
rect 149790 567196 149796 567248
rect 149848 567236 149854 567248
rect 151814 567236 151820 567248
rect 149848 567208 151820 567236
rect 149848 567196 149854 567208
rect 151814 567196 151820 567208
rect 151872 567196 151878 567248
rect 57054 566720 57060 566772
rect 57112 566760 57118 566772
rect 62114 566760 62120 566772
rect 57112 566732 62120 566760
rect 57112 566720 57118 566732
rect 62114 566720 62120 566732
rect 62172 566720 62178 566772
rect 156598 566720 156604 566772
rect 156656 566760 156662 566772
rect 213178 566760 213184 566772
rect 156656 566732 213184 566760
rect 156656 566720 156662 566732
rect 213178 566720 213184 566732
rect 213236 566720 213242 566772
rect 269114 566720 269120 566772
rect 269172 566760 269178 566772
rect 317138 566760 317144 566772
rect 269172 566732 317144 566760
rect 269172 566720 269178 566732
rect 317138 566720 317144 566732
rect 317196 566720 317202 566772
rect 125686 566652 125692 566704
rect 125744 566692 125750 566704
rect 211430 566692 211436 566704
rect 125744 566664 211436 566692
rect 125744 566652 125750 566664
rect 211430 566652 211436 566664
rect 211488 566652 211494 566704
rect 227714 566652 227720 566704
rect 227772 566692 227778 566704
rect 300946 566692 300952 566704
rect 227772 566664 300952 566692
rect 227772 566652 227778 566664
rect 300946 566652 300952 566664
rect 301004 566652 301010 566704
rect 57514 566584 57520 566636
rect 57572 566624 57578 566636
rect 82906 566624 82912 566636
rect 57572 566596 82912 566624
rect 57572 566584 57578 566596
rect 82906 566584 82912 566596
rect 82964 566584 82970 566636
rect 84194 566584 84200 566636
rect 84252 566624 84258 566636
rect 122098 566624 122104 566636
rect 84252 566596 122104 566624
rect 84252 566584 84258 566596
rect 122098 566584 122104 566596
rect 122156 566584 122162 566636
rect 200114 566584 200120 566636
rect 200172 566624 200178 566636
rect 302234 566624 302240 566636
rect 200172 566596 302240 566624
rect 200172 566584 200178 566596
rect 302234 566584 302240 566596
rect 302292 566584 302298 566636
rect 58526 566516 58532 566568
rect 58584 566556 58590 566568
rect 110414 566556 110420 566568
rect 58584 566528 110420 566556
rect 58584 566516 58590 566528
rect 110414 566516 110420 566528
rect 110472 566516 110478 566568
rect 180978 566516 180984 566568
rect 181036 566556 181042 566568
rect 301406 566556 301412 566568
rect 181036 566528 301412 566556
rect 181036 566516 181042 566528
rect 301406 566516 301412 566528
rect 301464 566516 301470 566568
rect 64874 566448 64880 566500
rect 64932 566488 64938 566500
rect 122006 566488 122012 566500
rect 64932 566460 122012 566488
rect 64932 566448 64938 566460
rect 122006 566448 122012 566460
rect 122064 566448 122070 566500
rect 148502 566448 148508 566500
rect 148560 566488 148566 566500
rect 160186 566488 160192 566500
rect 148560 566460 160192 566488
rect 148560 566448 148566 566460
rect 160186 566448 160192 566460
rect 160244 566448 160250 566500
rect 179506 566448 179512 566500
rect 179564 566488 179570 566500
rect 301590 566488 301596 566500
rect 179564 566460 301596 566488
rect 179564 566448 179570 566460
rect 301590 566448 301596 566460
rect 301648 566448 301654 566500
rect 148686 565836 148692 565888
rect 148744 565876 148750 565888
rect 150526 565876 150532 565888
rect 148744 565848 150532 565876
rect 148744 565836 148750 565848
rect 150526 565836 150532 565848
rect 150584 565836 150590 565888
rect 161566 565564 161572 565616
rect 161624 565604 161630 565616
rect 178034 565604 178040 565616
rect 161624 565576 178040 565604
rect 161624 565564 161630 565576
rect 178034 565564 178040 565576
rect 178092 565564 178098 565616
rect 82722 565496 82728 565548
rect 82780 565536 82786 565548
rect 89714 565536 89720 565548
rect 82780 565508 89720 565536
rect 82780 565496 82786 565508
rect 89714 565496 89720 565508
rect 89772 565496 89778 565548
rect 163038 565496 163044 565548
rect 163096 565536 163102 565548
rect 183830 565536 183836 565548
rect 163096 565508 183836 565536
rect 163096 565496 163102 565508
rect 183830 565496 183836 565508
rect 183888 565496 183894 565548
rect 235442 565496 235448 565548
rect 235500 565536 235506 565548
rect 248506 565536 248512 565548
rect 235500 565508 248512 565536
rect 235500 565496 235506 565508
rect 248506 565496 248512 565508
rect 248564 565496 248570 565548
rect 249058 565496 249064 565548
rect 249116 565536 249122 565548
rect 271230 565536 271236 565548
rect 249116 565508 271236 565536
rect 249116 565496 249122 565508
rect 271230 565496 271236 565508
rect 271288 565496 271294 565548
rect 74626 565428 74632 565480
rect 74684 565468 74690 565480
rect 96982 565468 96988 565480
rect 74684 565440 96988 565468
rect 74684 565428 74690 565440
rect 96982 565428 96988 565440
rect 97040 565428 97046 565480
rect 100202 565428 100208 565480
rect 100260 565468 100266 565480
rect 115198 565468 115204 565480
rect 100260 565440 115204 565468
rect 100260 565428 100266 565440
rect 115198 565428 115204 565440
rect 115256 565428 115262 565480
rect 143534 565428 143540 565480
rect 143592 565468 143598 565480
rect 166442 565468 166448 565480
rect 143592 565440 166448 565468
rect 143592 565428 143598 565440
rect 166442 565428 166448 565440
rect 166500 565428 166506 565480
rect 173894 565428 173900 565480
rect 173952 565468 173958 565480
rect 189626 565468 189632 565480
rect 173952 565440 189632 565468
rect 173952 565428 173958 565440
rect 189626 565428 189632 565440
rect 189684 565428 189690 565480
rect 230474 565428 230480 565480
rect 230532 565468 230538 565480
rect 259638 565468 259644 565480
rect 230532 565440 259644 565468
rect 230532 565428 230538 565440
rect 259638 565428 259644 565440
rect 259696 565428 259702 565480
rect 269758 565428 269764 565480
rect 269816 565468 269822 565480
rect 282914 565468 282920 565480
rect 269816 565440 282920 565468
rect 269816 565428 269822 565440
rect 282914 565428 282920 565440
rect 282972 565428 282978 565480
rect 77018 565360 77024 565412
rect 77076 565400 77082 565412
rect 84838 565400 84844 565412
rect 77076 565372 84844 565400
rect 77076 565360 77082 565372
rect 84838 565360 84844 565372
rect 84896 565360 84902 565412
rect 86034 565360 86040 565412
rect 86092 565400 86098 565412
rect 108390 565400 108396 565412
rect 86092 565372 108396 565400
rect 86092 565360 86098 565372
rect 108390 565360 108396 565372
rect 108448 565360 108454 565412
rect 154666 565360 154672 565412
rect 154724 565400 154730 565412
rect 181254 565400 181260 565412
rect 154724 565372 181260 565400
rect 154724 565360 154730 565372
rect 181254 565360 181260 565372
rect 181312 565360 181318 565412
rect 187786 565360 187792 565412
rect 187844 565400 187850 565412
rect 198734 565400 198740 565412
rect 187844 565372 198740 565400
rect 187844 565360 187850 565372
rect 198734 565360 198740 565372
rect 198792 565360 198798 565412
rect 227806 565360 227812 565412
rect 227864 565400 227870 565412
rect 265526 565400 265532 565412
rect 227864 565372 265532 565400
rect 227864 565360 227870 565372
rect 265526 565360 265532 565372
rect 265584 565360 265590 565412
rect 273346 565360 273352 565412
rect 273404 565400 273410 565412
rect 296990 565400 296996 565412
rect 273404 565372 296996 565400
rect 273404 565360 273410 565372
rect 296990 565360 296996 565372
rect 297048 565360 297054 565412
rect 79870 565292 79876 565344
rect 79928 565332 79934 565344
rect 114646 565332 114652 565344
rect 79928 565304 114652 565332
rect 79928 565292 79934 565304
rect 114646 565292 114652 565304
rect 114704 565292 114710 565344
rect 158714 565292 158720 565344
rect 158772 565332 158778 565344
rect 192846 565332 192852 565344
rect 158772 565304 192852 565332
rect 158772 565292 158778 565304
rect 192846 565292 192852 565304
rect 192904 565292 192910 565344
rect 196618 565292 196624 565344
rect 196676 565332 196682 565344
rect 210234 565332 210240 565344
rect 196676 565304 210240 565332
rect 196676 565292 196682 565304
rect 210234 565292 210240 565304
rect 210292 565292 210298 565344
rect 231946 565292 231952 565344
rect 232004 565332 232010 565344
rect 279694 565332 279700 565344
rect 232004 565304 279700 565332
rect 232004 565292 232010 565304
rect 279694 565292 279700 565304
rect 279752 565292 279758 565344
rect 291838 565292 291844 565344
rect 291896 565332 291902 565344
rect 300302 565332 300308 565344
rect 291896 565304 300308 565332
rect 291896 565292 291902 565304
rect 300302 565292 300308 565304
rect 300360 565292 300366 565344
rect 71314 565224 71320 565276
rect 71372 565264 71378 565276
rect 109678 565264 109684 565276
rect 71372 565236 109684 565264
rect 71372 565224 71378 565236
rect 109678 565224 109684 565236
rect 109736 565224 109742 565276
rect 129734 565224 129740 565276
rect 129792 565264 129798 565276
rect 163866 565264 163872 565276
rect 129792 565236 163872 565264
rect 129792 565224 129798 565236
rect 163866 565224 163872 565236
rect 163924 565224 163930 565276
rect 184198 565224 184204 565276
rect 184256 565264 184262 565276
rect 213086 565264 213092 565276
rect 184256 565236 213092 565264
rect 184256 565224 184262 565236
rect 213086 565224 213092 565236
rect 213144 565224 213150 565276
rect 219434 565224 219440 565276
rect 219492 565264 219498 565276
rect 268102 565264 268108 565276
rect 219492 565236 268108 565264
rect 219492 565224 219498 565236
rect 268102 565224 268108 565236
rect 268160 565224 268166 565276
rect 269206 565224 269212 565276
rect 269264 565264 269270 565276
rect 307202 565264 307208 565276
rect 269264 565236 307208 565264
rect 269264 565224 269270 565236
rect 307202 565224 307208 565236
rect 307260 565224 307266 565276
rect 60274 565156 60280 565208
rect 60332 565196 60338 565208
rect 104158 565196 104164 565208
rect 60332 565168 104164 565196
rect 60332 565156 60338 565168
rect 104158 565156 104164 565168
rect 104216 565156 104222 565208
rect 112438 565156 112444 565208
rect 112496 565196 112502 565208
rect 117406 565196 117412 565208
rect 112496 565168 117412 565196
rect 112496 565156 112502 565168
rect 117406 565156 117412 565168
rect 117464 565156 117470 565208
rect 132586 565156 132592 565208
rect 132644 565196 132650 565208
rect 187050 565196 187056 565208
rect 132644 565168 187056 565196
rect 132644 565156 132650 565168
rect 187050 565156 187056 565168
rect 187108 565156 187114 565208
rect 195238 565156 195244 565208
rect 195296 565196 195302 565208
rect 212718 565196 212724 565208
rect 195296 565168 212724 565196
rect 195296 565156 195302 565168
rect 212718 565156 212724 565168
rect 212776 565156 212782 565208
rect 222286 565156 222292 565208
rect 222344 565196 222350 565208
rect 273806 565196 273812 565208
rect 222344 565168 273812 565196
rect 222344 565156 222350 565168
rect 273806 565156 273812 565168
rect 273864 565156 273870 565208
rect 280154 565156 280160 565208
rect 280212 565196 280218 565208
rect 322474 565196 322480 565208
rect 280212 565168 322480 565196
rect 280212 565156 280218 565168
rect 322474 565156 322480 565168
rect 322532 565156 322538 565208
rect 62850 565088 62856 565140
rect 62908 565128 62914 565140
rect 108298 565128 108304 565140
rect 62908 565100 108304 565128
rect 62908 565088 62914 565100
rect 108298 565088 108304 565100
rect 108356 565088 108362 565140
rect 110506 565088 110512 565140
rect 110564 565128 110570 565140
rect 120718 565128 120724 565140
rect 110564 565100 120724 565128
rect 110564 565088 110570 565100
rect 120718 565088 120724 565100
rect 120776 565088 120782 565140
rect 133966 565088 133972 565140
rect 134024 565128 134030 565140
rect 207014 565128 207020 565140
rect 134024 565100 207020 565128
rect 134024 565088 134030 565100
rect 207014 565088 207020 565100
rect 207072 565088 207078 565140
rect 220814 565088 220820 565140
rect 220872 565128 220878 565140
rect 239766 565128 239772 565140
rect 220872 565100 239772 565128
rect 220872 565088 220878 565100
rect 239766 565088 239772 565100
rect 239824 565088 239830 565140
rect 259454 565088 259460 565140
rect 259512 565128 259518 565140
rect 321094 565128 321100 565140
rect 259512 565100 321100 565128
rect 259512 565088 259518 565100
rect 321094 565088 321100 565100
rect 321152 565088 321158 565140
rect 94498 564884 94504 564936
rect 94556 564924 94562 564936
rect 102778 564924 102784 564936
rect 94556 564896 102784 564924
rect 94556 564884 94562 564896
rect 102778 564884 102784 564896
rect 102836 564884 102842 564936
rect 150342 564544 150348 564596
rect 150400 564584 150406 564596
rect 151170 564584 151176 564596
rect 150400 564556 151176 564584
rect 150400 564544 150406 564556
rect 151170 564544 151176 564556
rect 151228 564544 151234 564596
rect 216674 564544 216680 564596
rect 216732 564584 216738 564596
rect 220354 564584 220360 564596
rect 216732 564556 220360 564584
rect 216732 564544 216738 564556
rect 220354 564544 220360 564556
rect 220412 564544 220418 564596
rect 71774 564408 71780 564460
rect 71832 564448 71838 564460
rect 73798 564448 73804 564460
rect 71832 564420 73804 564448
rect 71832 564408 71838 564420
rect 73798 564408 73804 564420
rect 73856 564408 73862 564460
rect 100754 564408 100760 564460
rect 100812 564448 100818 564460
rect 102870 564448 102876 564460
rect 100812 564420 102876 564448
rect 100812 564408 100818 564420
rect 102870 564408 102876 564420
rect 102928 564408 102934 564460
rect 116578 564408 116584 564460
rect 116636 564448 116642 564460
rect 120166 564448 120172 564460
rect 116636 564420 120172 564448
rect 116636 564408 116642 564420
rect 120166 564408 120172 564420
rect 120224 564408 120230 564460
rect 191098 564408 191104 564460
rect 191156 564448 191162 564460
rect 195422 564448 195428 564460
rect 191156 564420 195428 564448
rect 191156 564408 191162 564420
rect 195422 564408 195428 564420
rect 195480 564408 195486 564460
rect 197998 564408 198004 564460
rect 198056 564448 198062 564460
rect 201494 564448 201500 564460
rect 198056 564420 201500 564448
rect 198056 564408 198062 564420
rect 201494 564408 201500 564420
rect 201552 564408 201558 564460
rect 202138 564408 202144 564460
rect 202196 564448 202202 564460
rect 204438 564448 204444 564460
rect 202196 564420 204444 564448
rect 202196 564408 202202 564420
rect 204438 564408 204444 564420
rect 204496 564408 204502 564460
rect 244918 564408 244924 564460
rect 244976 564448 244982 564460
rect 250622 564448 250628 564460
rect 244976 564420 250628 564448
rect 244976 564408 244982 564420
rect 250622 564408 250628 564420
rect 250680 564408 250686 564460
rect 282178 564408 282184 564460
rect 282236 564448 282242 564460
rect 288710 564448 288716 564460
rect 282236 564420 288716 564448
rect 282236 564408 282242 564420
rect 288710 564408 288716 564420
rect 288768 564408 288774 564460
rect 200206 563932 200212 563984
rect 200264 563972 200270 563984
rect 239582 563972 239588 563984
rect 200264 563944 239588 563972
rect 200264 563932 200270 563944
rect 239582 563932 239588 563944
rect 239640 563932 239646 563984
rect 191834 563864 191840 563916
rect 191892 563904 191898 563916
rect 238846 563904 238852 563916
rect 191892 563876 238852 563904
rect 191892 563864 191898 563876
rect 238846 563864 238852 563876
rect 238904 563864 238910 563916
rect 263594 563864 263600 563916
rect 263652 563904 263658 563916
rect 322382 563904 322388 563916
rect 263652 563876 322388 563904
rect 263652 563864 263658 563876
rect 322382 563864 322388 563876
rect 322440 563864 322446 563916
rect 58894 563796 58900 563848
rect 58952 563836 58958 563848
rect 91186 563836 91192 563848
rect 58952 563808 91192 563836
rect 58952 563796 58958 563808
rect 91186 563796 91192 563808
rect 91244 563796 91250 563848
rect 126974 563796 126980 563848
rect 127032 563836 127038 563848
rect 211798 563836 211804 563848
rect 127032 563808 211804 563836
rect 127032 563796 127038 563808
rect 211798 563796 211804 563808
rect 211856 563796 211862 563848
rect 215386 563796 215392 563848
rect 215444 563836 215450 563848
rect 301498 563836 301504 563848
rect 215444 563808 301504 563836
rect 215444 563796 215450 563808
rect 301498 563796 301504 563808
rect 301556 563796 301562 563848
rect 69014 563728 69020 563780
rect 69072 563768 69078 563780
rect 123386 563768 123392 563780
rect 69072 563740 123392 563768
rect 69072 563728 69078 563740
rect 123386 563728 123392 563740
rect 123444 563728 123450 563780
rect 146846 563728 146852 563780
rect 146904 563768 146910 563780
rect 165614 563768 165620 563780
rect 146904 563740 165620 563768
rect 146904 563728 146910 563740
rect 165614 563728 165620 563740
rect 165672 563728 165678 563780
rect 180886 563728 180892 563780
rect 180944 563768 180950 563780
rect 301222 563768 301228 563780
rect 180944 563740 301228 563768
rect 180944 563728 180950 563740
rect 301222 563728 301228 563740
rect 301280 563728 301286 563780
rect 10318 563660 10324 563712
rect 10376 563700 10382 563712
rect 321554 563700 321560 563712
rect 10376 563672 321560 563700
rect 10376 563660 10382 563672
rect 321554 563660 321560 563672
rect 321612 563660 321618 563712
rect 273254 562640 273260 562692
rect 273312 562680 273318 562692
rect 322290 562680 322296 562692
rect 273312 562652 322296 562680
rect 273312 562640 273318 562652
rect 322290 562640 322296 562652
rect 322348 562640 322354 562692
rect 204254 562572 204260 562624
rect 204312 562612 204318 562624
rect 239490 562612 239496 562624
rect 204312 562584 239496 562612
rect 204312 562572 204318 562584
rect 239490 562572 239496 562584
rect 239548 562572 239554 562624
rect 255314 562572 255320 562624
rect 255372 562612 255378 562624
rect 324774 562612 324780 562624
rect 255372 562584 324780 562612
rect 255372 562572 255378 562584
rect 324774 562572 324780 562584
rect 324832 562572 324838 562624
rect 157518 562504 157524 562556
rect 157576 562544 157582 562556
rect 212534 562544 212540 562556
rect 157576 562516 212540 562544
rect 157576 562504 157582 562516
rect 212534 562504 212540 562516
rect 212592 562504 212598 562556
rect 242894 562504 242900 562556
rect 242952 562544 242958 562556
rect 318058 562544 318064 562556
rect 242952 562516 318064 562544
rect 242952 562504 242958 562516
rect 318058 562504 318064 562516
rect 318116 562504 318122 562556
rect 68738 562436 68744 562488
rect 68796 562476 68802 562488
rect 106918 562476 106924 562488
rect 68796 562448 106924 562476
rect 68796 562436 68802 562448
rect 106918 562436 106924 562448
rect 106976 562436 106982 562488
rect 111886 562436 111892 562488
rect 111944 562476 111950 562488
rect 123018 562476 123024 562488
rect 111944 562448 123024 562476
rect 111944 562436 111950 562448
rect 123018 562436 123024 562448
rect 123076 562436 123082 562488
rect 191926 562436 191932 562488
rect 191984 562476 191990 562488
rect 273346 562476 273352 562488
rect 191984 562448 273352 562476
rect 191984 562436 191990 562448
rect 273346 562436 273352 562448
rect 273404 562436 273410 562488
rect 59446 562368 59452 562420
rect 59504 562408 59510 562420
rect 75914 562408 75920 562420
rect 59504 562380 75920 562408
rect 59504 562368 59510 562380
rect 75914 562368 75920 562380
rect 75972 562368 75978 562420
rect 78766 562368 78772 562420
rect 78824 562408 78830 562420
rect 121178 562408 121184 562420
rect 78824 562380 121184 562408
rect 78824 562368 78830 562380
rect 121178 562368 121184 562380
rect 121236 562368 121242 562420
rect 184934 562368 184940 562420
rect 184992 562408 184998 562420
rect 294414 562408 294420 562420
rect 184992 562380 294420 562408
rect 184992 562368 184998 562380
rect 294414 562368 294420 562380
rect 294472 562368 294478 562420
rect 69106 562300 69112 562352
rect 69164 562340 69170 562352
rect 114554 562340 114560 562352
rect 69164 562312 114560 562340
rect 69164 562300 69170 562312
rect 114554 562300 114560 562312
rect 114612 562300 114618 562352
rect 118694 562300 118700 562352
rect 118752 562340 118758 562352
rect 154850 562340 154856 562352
rect 118752 562312 154856 562340
rect 118752 562300 118758 562312
rect 154850 562300 154856 562312
rect 154908 562300 154914 562352
rect 186314 562300 186320 562352
rect 186372 562340 186378 562352
rect 302786 562340 302792 562352
rect 186372 562312 302792 562340
rect 186372 562300 186378 562312
rect 302786 562300 302792 562312
rect 302844 562300 302850 562352
rect 198734 561212 198740 561264
rect 198792 561252 198798 561264
rect 239398 561252 239404 561264
rect 198792 561224 239404 561252
rect 198792 561212 198798 561224
rect 239398 561212 239404 561224
rect 239456 561212 239462 561264
rect 266446 561212 266452 561264
rect 266504 561252 266510 561264
rect 307018 561252 307024 561264
rect 266504 561224 307024 561252
rect 266504 561212 266510 561224
rect 307018 561212 307024 561224
rect 307076 561212 307082 561264
rect 148226 561144 148232 561196
rect 148284 561184 148290 561196
rect 158806 561184 158812 561196
rect 148284 561156 158812 561184
rect 148284 561144 148290 561156
rect 158806 561144 158812 561156
rect 158864 561144 158870 561196
rect 176654 561144 176660 561196
rect 176712 561184 176718 561196
rect 217502 561184 217508 561196
rect 176712 561156 217508 561184
rect 176712 561144 176718 561156
rect 217502 561144 217508 561156
rect 217560 561144 217566 561196
rect 251174 561144 251180 561196
rect 251232 561184 251238 561196
rect 323946 561184 323952 561196
rect 251232 561156 323952 561184
rect 251232 561144 251238 561156
rect 323946 561144 323952 561156
rect 324004 561144 324010 561196
rect 59262 561076 59268 561128
rect 59320 561116 59326 561128
rect 92566 561116 92572 561128
rect 59320 561088 92572 561116
rect 59320 561076 59326 561088
rect 92566 561076 92572 561088
rect 92624 561076 92630 561128
rect 138014 561076 138020 561128
rect 138072 561116 138078 561128
rect 211614 561116 211620 561128
rect 138072 561088 211620 561116
rect 138072 561076 138078 561088
rect 211614 561076 211620 561088
rect 211672 561076 211678 561128
rect 240134 561076 240140 561128
rect 240192 561116 240198 561128
rect 313918 561116 313924 561128
rect 240192 561088 313924 561116
rect 240192 561076 240198 561088
rect 313918 561076 313924 561088
rect 313976 561076 313982 561128
rect 70394 561008 70400 561060
rect 70452 561048 70458 561060
rect 121914 561048 121920 561060
rect 70452 561020 121920 561048
rect 70452 561008 70458 561020
rect 121914 561008 121920 561020
rect 121972 561008 121978 561060
rect 147030 561008 147036 561060
rect 147088 561048 147094 561060
rect 168374 561048 168380 561060
rect 147088 561020 168380 561048
rect 147088 561008 147094 561020
rect 168374 561008 168380 561020
rect 168432 561008 168438 561060
rect 187694 561008 187700 561060
rect 187752 561048 187758 561060
rect 301038 561048 301044 561060
rect 187752 561020 301044 561048
rect 187752 561008 187758 561020
rect 301038 561008 301044 561020
rect 301096 561008 301102 561060
rect 63586 560940 63592 560992
rect 63644 560980 63650 560992
rect 122834 560980 122840 560992
rect 63644 560952 122840 560980
rect 63644 560940 63650 560952
rect 122834 560940 122840 560952
rect 122892 560940 122898 560992
rect 147306 560940 147312 560992
rect 147364 560980 147370 560992
rect 175366 560980 175372 560992
rect 147364 560952 175372 560980
rect 147364 560940 147370 560952
rect 175366 560940 175372 560952
rect 175424 560940 175430 560992
rect 182174 560940 182180 560992
rect 182232 560980 182238 560992
rect 301682 560980 301688 560992
rect 182232 560952 301688 560980
rect 182232 560940 182238 560952
rect 301682 560940 301688 560952
rect 301740 560940 301746 560992
rect 201494 559784 201500 559836
rect 201552 559824 201558 559836
rect 256694 559824 256700 559836
rect 201552 559796 256700 559824
rect 201552 559784 201558 559796
rect 256694 559784 256700 559796
rect 256752 559784 256758 559836
rect 88426 559716 88432 559768
rect 88484 559756 88490 559768
rect 103514 559756 103520 559768
rect 88484 559728 103520 559756
rect 88484 559716 88490 559728
rect 103514 559716 103520 559728
rect 103572 559716 103578 559768
rect 176746 559716 176752 559768
rect 176804 559756 176810 559768
rect 244274 559756 244280 559768
rect 176804 559728 244280 559756
rect 176804 559716 176810 559728
rect 244274 559716 244280 559728
rect 244332 559716 244338 559768
rect 57238 559648 57244 559700
rect 57296 559688 57302 559700
rect 89806 559688 89812 559700
rect 57296 559660 89812 559688
rect 57296 559648 57302 559660
rect 89806 559648 89812 559660
rect 89864 559648 89870 559700
rect 190454 559648 190460 559700
rect 190512 559688 190518 559700
rect 277486 559688 277492 559700
rect 190512 559660 277492 559688
rect 190512 559648 190518 559660
rect 277486 559648 277492 559660
rect 277544 559648 277550 559700
rect 85666 559580 85672 559632
rect 85724 559620 85730 559632
rect 121822 559620 121828 559632
rect 85724 559592 121828 559620
rect 85724 559580 85730 559592
rect 121822 559580 121828 559592
rect 121880 559580 121886 559632
rect 122834 559580 122840 559632
rect 122892 559620 122898 559632
rect 211338 559620 211344 559632
rect 122892 559592 211344 559620
rect 122892 559580 122898 559592
rect 211338 559580 211344 559592
rect 211396 559580 211402 559632
rect 244274 559580 244280 559632
rect 244332 559620 244338 559632
rect 319438 559620 319444 559632
rect 244332 559592 319444 559620
rect 244332 559580 244338 559592
rect 319438 559580 319444 559592
rect 319496 559580 319502 559632
rect 65058 559512 65064 559564
rect 65116 559552 65122 559564
rect 123110 559552 123116 559564
rect 65116 559524 123116 559552
rect 65116 559512 65122 559524
rect 123110 559512 123116 559524
rect 123168 559512 123174 559564
rect 149054 559512 149060 559564
rect 149112 559552 149118 559564
rect 160278 559552 160284 559564
rect 149112 559524 160284 559552
rect 149112 559512 149118 559524
rect 160278 559512 160284 559524
rect 160336 559512 160342 559564
rect 195974 559512 195980 559564
rect 196032 559552 196038 559564
rect 302602 559552 302608 559564
rect 196032 559524 302608 559552
rect 196032 559512 196038 559524
rect 302602 559512 302608 559524
rect 302660 559512 302666 559564
rect 267734 558900 267740 558952
rect 267792 558940 267798 558952
rect 321554 558940 321560 558952
rect 267792 558912 321560 558940
rect 267792 558900 267798 558912
rect 321554 558900 321560 558912
rect 321612 558900 321618 558952
rect 190546 558424 190552 558476
rect 190604 558464 190610 558476
rect 222838 558464 222844 558476
rect 190604 558436 222844 558464
rect 190604 558424 190610 558436
rect 222838 558424 222844 558436
rect 222896 558424 222902 558476
rect 270494 558424 270500 558476
rect 270552 558464 270558 558476
rect 309778 558464 309784 558476
rect 270552 558436 309784 558464
rect 270552 558424 270558 558436
rect 309778 558424 309784 558436
rect 309836 558424 309842 558476
rect 88426 558356 88432 558408
rect 88484 558396 88490 558408
rect 104894 558396 104900 558408
rect 88484 558368 104900 558396
rect 88484 558356 88490 558368
rect 104894 558356 104900 558368
rect 104952 558356 104958 558408
rect 178034 558356 178040 558408
rect 178092 558396 178098 558408
rect 236730 558396 236736 558408
rect 178092 558368 236736 558396
rect 178092 558356 178098 558368
rect 236730 558356 236736 558368
rect 236788 558356 236794 558408
rect 249794 558356 249800 558408
rect 249852 558396 249858 558408
rect 307110 558396 307116 558408
rect 249852 558368 307116 558396
rect 249852 558356 249858 558368
rect 307110 558356 307116 558368
rect 307168 558356 307174 558408
rect 98638 558288 98644 558340
rect 98696 558328 98702 558340
rect 123294 558328 123300 558340
rect 98696 558300 123300 558328
rect 98696 558288 98702 558300
rect 123294 558288 123300 558300
rect 123352 558288 123358 558340
rect 205634 558288 205640 558340
rect 205692 558328 205698 558340
rect 285674 558328 285680 558340
rect 205692 558300 285680 558328
rect 205692 558288 205698 558300
rect 285674 558288 285680 558300
rect 285732 558288 285738 558340
rect 80054 558220 80060 558272
rect 80112 558260 80118 558272
rect 120810 558260 120816 558272
rect 80112 558232 120816 558260
rect 80112 558220 80118 558232
rect 120810 558220 120816 558232
rect 120868 558220 120874 558272
rect 122926 558220 122932 558272
rect 122984 558260 122990 558272
rect 211706 558260 211712 558272
rect 122984 558232 211712 558260
rect 122984 558220 122990 558232
rect 211706 558220 211712 558232
rect 211764 558220 211770 558272
rect 252554 558220 252560 558272
rect 252612 558260 252618 558272
rect 323854 558260 323860 558272
rect 252612 558232 323860 558260
rect 252612 558220 252618 558232
rect 323854 558220 323860 558232
rect 323912 558220 323918 558272
rect 59538 558152 59544 558204
rect 59596 558192 59602 558204
rect 100846 558192 100852 558204
rect 59596 558164 100852 558192
rect 59596 558152 59602 558164
rect 100846 558152 100852 558164
rect 100904 558152 100910 558204
rect 131114 558152 131120 558204
rect 131172 558192 131178 558204
rect 187786 558192 187792 558204
rect 131172 558164 187792 558192
rect 131172 558152 131178 558164
rect 187786 558152 187792 558164
rect 187844 558152 187850 558204
rect 196066 558152 196072 558204
rect 196124 558192 196130 558204
rect 302970 558192 302976 558204
rect 196124 558164 302976 558192
rect 196124 558152 196130 558164
rect 302970 558152 302976 558164
rect 303028 558152 303034 558204
rect 199194 557064 199200 557116
rect 199252 557104 199258 557116
rect 232498 557104 232504 557116
rect 199252 557076 232504 557104
rect 199252 557064 199258 557076
rect 232498 557064 232504 557076
rect 232556 557064 232562 557116
rect 80974 556996 80980 557048
rect 81032 557036 81038 557048
rect 121086 557036 121092 557048
rect 81032 557008 121092 557036
rect 81032 556996 81038 557008
rect 121086 556996 121092 557008
rect 121144 556996 121150 557048
rect 189902 556996 189908 557048
rect 189960 557036 189966 557048
rect 238202 557036 238208 557048
rect 189960 557008 238208 557036
rect 189960 556996 189966 557008
rect 238202 556996 238208 557008
rect 238260 556996 238266 557048
rect 57422 556928 57428 556980
rect 57480 556968 57486 556980
rect 81710 556968 81716 556980
rect 57480 556940 81716 556968
rect 57480 556928 57486 556940
rect 81710 556928 81716 556940
rect 81768 556928 81774 556980
rect 137186 556928 137192 556980
rect 137244 556968 137250 556980
rect 212810 556968 212816 556980
rect 137244 556940 212816 556968
rect 137244 556928 137250 556940
rect 212810 556928 212816 556940
rect 212868 556928 212874 556980
rect 250806 556928 250812 556980
rect 250864 556968 250870 556980
rect 323762 556968 323768 556980
rect 250864 556940 323768 556968
rect 250864 556928 250870 556940
rect 323762 556928 323768 556940
rect 323820 556928 323826 556980
rect 121086 556860 121092 556912
rect 121144 556900 121150 556912
rect 197998 556900 198004 556912
rect 121144 556872 198004 556900
rect 121144 556860 121150 556872
rect 197998 556860 198004 556872
rect 198056 556860 198062 556912
rect 202230 556860 202236 556912
rect 202288 556900 202294 556912
rect 302878 556900 302884 556912
rect 202288 556872 302884 556900
rect 202288 556860 202294 556872
rect 302878 556860 302884 556872
rect 302936 556860 302942 556912
rect 59078 556792 59084 556844
rect 59136 556832 59142 556844
rect 102502 556832 102508 556844
rect 59136 556804 102508 556832
rect 59136 556792 59142 556804
rect 102502 556792 102508 556804
rect 102560 556792 102566 556844
rect 147214 556792 147220 556844
rect 147272 556832 147278 556844
rect 174906 556832 174912 556844
rect 147272 556804 174912 556832
rect 147272 556792 147278 556804
rect 174906 556792 174912 556804
rect 174964 556792 174970 556844
rect 179138 556792 179144 556844
rect 179196 556832 179202 556844
rect 291286 556832 291292 556844
rect 179196 556804 291292 556832
rect 179196 556792 179202 556804
rect 291286 556792 291292 556804
rect 291344 556792 291350 556844
rect 125594 555772 125600 555824
rect 125652 555812 125658 555824
rect 126882 555812 126888 555824
rect 125652 555784 126888 555812
rect 125652 555772 125658 555784
rect 126882 555772 126888 555784
rect 126940 555772 126946 555824
rect 197814 555636 197820 555688
rect 197872 555676 197878 555688
rect 216030 555676 216036 555688
rect 197872 555648 216036 555676
rect 197872 555636 197878 555648
rect 216030 555636 216036 555648
rect 216088 555636 216094 555688
rect 73154 555568 73160 555620
rect 73212 555608 73218 555620
rect 107654 555608 107660 555620
rect 73212 555580 107660 555608
rect 73212 555568 73218 555580
rect 107654 555568 107660 555580
rect 107712 555568 107718 555620
rect 142614 555568 142620 555620
rect 142672 555608 142678 555620
rect 212994 555608 213000 555620
rect 142672 555580 213000 555608
rect 142672 555568 142678 555580
rect 212994 555568 213000 555580
rect 213052 555568 213058 555620
rect 282362 555568 282368 555620
rect 282420 555608 282426 555620
rect 305730 555608 305736 555620
rect 282420 555580 305736 555608
rect 282420 555568 282426 555580
rect 305730 555568 305736 555580
rect 305788 555568 305794 555620
rect 189166 555500 189172 555552
rect 189224 555540 189230 555552
rect 282178 555540 282184 555552
rect 189224 555512 282184 555540
rect 189224 555500 189230 555512
rect 282178 555500 282184 555512
rect 282236 555500 282242 555552
rect 283742 555500 283748 555552
rect 283800 555540 283806 555552
rect 312630 555540 312636 555552
rect 283800 555512 312636 555540
rect 283800 555500 283806 555512
rect 312630 555500 312636 555512
rect 312688 555500 312694 555552
rect 59170 555432 59176 555484
rect 59228 555472 59234 555484
rect 108206 555472 108212 555484
rect 59228 555444 108212 555472
rect 59228 555432 59234 555444
rect 108206 555432 108212 555444
rect 108264 555432 108270 555484
rect 187050 555432 187056 555484
rect 187108 555472 187114 555484
rect 302418 555472 302424 555484
rect 187108 555444 302424 555472
rect 187108 555432 187114 555444
rect 302418 555432 302424 555444
rect 302476 555432 302482 555484
rect 21358 554752 21364 554804
rect 21416 554792 21422 554804
rect 321554 554792 321560 554804
rect 21416 554764 321560 554792
rect 21416 554752 21422 554764
rect 321554 554752 321560 554764
rect 321612 554752 321618 554804
rect 193490 554344 193496 554396
rect 193548 554384 193554 554396
rect 217410 554384 217416 554396
rect 193548 554356 217416 554384
rect 193548 554344 193554 554356
rect 217410 554344 217416 554356
rect 217468 554344 217474 554396
rect 206370 554276 206376 554328
rect 206428 554316 206434 554328
rect 262214 554316 262220 554328
rect 206428 554288 262220 554316
rect 206428 554276 206434 554288
rect 262214 554276 262220 554288
rect 262272 554276 262278 554328
rect 279510 554276 279516 554328
rect 279568 554316 279574 554328
rect 311158 554316 311164 554328
rect 279568 554288 311164 554316
rect 279568 554276 279574 554288
rect 311158 554276 311164 554288
rect 311216 554276 311222 554328
rect 168374 554208 168380 554260
rect 168432 554248 168438 554260
rect 210694 554248 210700 554260
rect 168432 554220 210700 554248
rect 168432 554208 168438 554220
rect 210694 554208 210700 554220
rect 210752 554208 210758 554260
rect 257982 554208 257988 554260
rect 258040 554248 258046 554260
rect 321002 554248 321008 554260
rect 258040 554220 321008 554248
rect 258040 554208 258046 554220
rect 321002 554208 321008 554220
rect 321060 554208 321066 554260
rect 57790 554140 57796 554192
rect 57848 554180 57854 554192
rect 103238 554180 103244 554192
rect 57848 554152 103244 554180
rect 57848 554140 57854 554152
rect 103238 554140 103244 554152
rect 103296 554140 103302 554192
rect 151170 554140 151176 554192
rect 151228 554180 151234 554192
rect 163406 554180 163412 554192
rect 151228 554152 163412 554180
rect 151228 554140 151234 554152
rect 163406 554140 163412 554152
rect 163464 554140 163470 554192
rect 184934 554140 184940 554192
rect 184992 554180 184998 554192
rect 235350 554180 235356 554192
rect 184992 554152 235356 554180
rect 184992 554140 184998 554152
rect 235350 554140 235356 554152
rect 235408 554140 235414 554192
rect 246482 554140 246488 554192
rect 246540 554180 246546 554192
rect 312538 554180 312544 554192
rect 246540 554152 312544 554180
rect 246540 554140 246546 554152
rect 312538 554140 312544 554152
rect 312596 554140 312602 554192
rect 63126 554072 63132 554124
rect 63184 554112 63190 554124
rect 110598 554112 110604 554124
rect 63184 554084 110604 554112
rect 63184 554072 63190 554084
rect 110598 554072 110604 554084
rect 110656 554072 110662 554124
rect 127618 554072 127624 554124
rect 127676 554112 127682 554124
rect 202138 554112 202144 554124
rect 127676 554084 202144 554112
rect 127676 554072 127682 554084
rect 202138 554072 202144 554084
rect 202196 554072 202202 554124
rect 229278 554072 229284 554124
rect 229336 554112 229342 554124
rect 303062 554112 303068 554124
rect 229336 554084 303068 554112
rect 229336 554072 229342 554084
rect 303062 554072 303068 554084
rect 303120 554072 303126 554124
rect 71682 554004 71688 554056
rect 71740 554044 71746 554056
rect 121730 554044 121736 554056
rect 71740 554016 121736 554044
rect 71740 554004 71746 554016
rect 121730 554004 121736 554016
rect 121788 554004 121794 554056
rect 140498 554004 140504 554056
rect 140556 554044 140562 554056
rect 196618 554044 196624 554056
rect 140556 554016 196624 554044
rect 140556 554004 140562 554016
rect 196618 554004 196624 554016
rect 196676 554004 196682 554056
rect 198550 554004 198556 554056
rect 198608 554044 198614 554056
rect 291838 554044 291844 554056
rect 198608 554016 291844 554044
rect 198608 554004 198614 554016
rect 291838 554004 291844 554016
rect 291896 554004 291902 554056
rect 200206 553052 200212 553104
rect 200264 553092 200270 553104
rect 201402 553092 201408 553104
rect 200264 553064 201408 553092
rect 200264 553052 200270 553064
rect 201402 553052 201408 553064
rect 201460 553052 201466 553104
rect 210786 553024 210792 553036
rect 121840 552996 210792 553024
rect 103486 552928 113174 552956
rect 89806 552848 89812 552900
rect 89864 552888 89870 552900
rect 91002 552888 91008 552900
rect 89864 552860 91008 552888
rect 89864 552848 89870 552860
rect 91002 552848 91008 552860
rect 91060 552848 91066 552900
rect 88426 552780 88432 552832
rect 88484 552820 88490 552832
rect 89622 552820 89628 552832
rect 88484 552792 89628 552820
rect 88484 552780 88490 552792
rect 89622 552780 89628 552792
rect 89680 552780 89686 552832
rect 100754 552780 100760 552832
rect 100812 552820 100818 552832
rect 101766 552820 101772 552832
rect 100812 552792 101772 552820
rect 100812 552780 100818 552792
rect 101766 552780 101772 552792
rect 101824 552780 101830 552832
rect 67634 552712 67640 552764
rect 67692 552752 67698 552764
rect 68830 552752 68836 552764
rect 67692 552724 68836 552752
rect 67692 552712 67698 552724
rect 68830 552712 68836 552724
rect 68888 552712 68894 552764
rect 69014 552712 69020 552764
rect 69072 552752 69078 552764
rect 70302 552752 70308 552764
rect 69072 552724 70308 552752
rect 69072 552712 69078 552724
rect 70302 552712 70308 552724
rect 70360 552712 70366 552764
rect 78674 552712 78680 552764
rect 78732 552752 78738 552764
rect 79594 552752 79600 552764
rect 78732 552724 79600 552752
rect 78732 552712 78738 552724
rect 79594 552712 79600 552724
rect 79652 552712 79658 552764
rect 82446 552712 82452 552764
rect 82504 552752 82510 552764
rect 103486 552752 103514 552928
rect 112438 552888 112444 552900
rect 82504 552724 103514 552752
rect 103624 552860 112444 552888
rect 82504 552712 82510 552724
rect 76742 552644 76748 552696
rect 76800 552684 76806 552696
rect 103624 552684 103652 552860
rect 112438 552848 112444 552860
rect 112496 552848 112502 552900
rect 113146 552752 113174 552928
rect 116578 552752 116584 552764
rect 113146 552724 116584 552752
rect 116578 552712 116584 552724
rect 116636 552712 116642 552764
rect 121840 552696 121868 552996
rect 210786 552984 210792 552996
rect 210844 552984 210850 553036
rect 213546 552984 213552 553036
rect 213604 553024 213610 553036
rect 235258 553024 235264 553036
rect 213604 552996 235264 553024
rect 213604 552984 213610 552996
rect 235258 552984 235264 552996
rect 235316 552984 235322 553036
rect 173802 552916 173808 552968
rect 173860 552956 173866 552968
rect 213362 552956 213368 552968
rect 173860 552928 213368 552956
rect 173860 552916 173866 552928
rect 213362 552916 213368 552928
rect 213420 552916 213426 552968
rect 260098 552916 260104 552968
rect 260156 552956 260162 552968
rect 311250 552956 311256 552968
rect 260156 552928 311256 552956
rect 260156 552916 260162 552928
rect 311250 552916 311256 552928
rect 311308 552916 311314 552968
rect 211154 552888 211160 552900
rect 129752 552860 211160 552888
rect 122834 552712 122840 552764
rect 122892 552752 122898 552764
rect 124030 552752 124036 552764
rect 122892 552724 124036 552752
rect 122892 552712 122898 552724
rect 124030 552712 124036 552724
rect 124088 552712 124094 552764
rect 124214 552712 124220 552764
rect 124272 552752 124278 552764
rect 125410 552752 125416 552764
rect 124272 552724 125416 552752
rect 124272 552712 124278 552724
rect 125410 552712 125416 552724
rect 125468 552712 125474 552764
rect 126974 552712 126980 552764
rect 127032 552752 127038 552764
rect 128262 552752 128268 552764
rect 127032 552724 128268 552752
rect 127032 552712 127038 552724
rect 128262 552712 128268 552724
rect 128320 552712 128326 552764
rect 129752 552696 129780 552860
rect 211154 552848 211160 552860
rect 211212 552848 211218 552900
rect 217870 552848 217876 552900
rect 217928 552888 217934 552900
rect 269758 552888 269764 552900
rect 217928 552860 269764 552888
rect 217928 552848 217934 552860
rect 269758 552848 269764 552860
rect 269816 552848 269822 552900
rect 275186 552848 275192 552900
rect 275244 552888 275250 552900
rect 316770 552888 316776 552900
rect 275244 552860 316776 552888
rect 275244 552848 275250 552860
rect 316770 552848 316776 552860
rect 316828 552848 316834 552900
rect 146294 552780 146300 552832
rect 146352 552820 146358 552832
rect 213270 552820 213276 552832
rect 146352 552792 213276 552820
rect 146352 552780 146358 552792
rect 213270 552780 213276 552792
rect 213328 552780 213334 552832
rect 219434 552780 219440 552832
rect 219492 552820 219498 552832
rect 220722 552820 220728 552832
rect 219492 552792 220728 552820
rect 219492 552780 219498 552792
rect 220722 552780 220728 552792
rect 220780 552780 220786 552832
rect 222194 552780 222200 552832
rect 222252 552820 222258 552832
rect 222838 552820 222844 552832
rect 222252 552792 222844 552820
rect 222252 552780 222258 552792
rect 222838 552780 222844 552792
rect 222896 552780 222902 552832
rect 227714 552780 227720 552832
rect 227772 552820 227778 552832
rect 228634 552820 228640 552832
rect 227772 552792 228640 552820
rect 227772 552780 227778 552792
rect 228634 552780 228640 552792
rect 228692 552780 228698 552832
rect 231854 552780 231860 552832
rect 231912 552820 231918 552832
rect 232866 552820 232872 552832
rect 231912 552792 232872 552820
rect 231912 552780 231918 552792
rect 232866 552780 232872 552792
rect 232924 552780 232930 552832
rect 247954 552780 247960 552832
rect 248012 552820 248018 552832
rect 324866 552820 324872 552832
rect 248012 552792 324872 552820
rect 248012 552780 248018 552792
rect 324866 552780 324872 552792
rect 324924 552780 324930 552832
rect 140774 552712 140780 552764
rect 140832 552752 140838 552764
rect 141878 552752 141884 552764
rect 140832 552724 141884 552752
rect 140832 552712 140838 552724
rect 141878 552712 141884 552724
rect 141936 552712 141942 552764
rect 142154 552712 142160 552764
rect 142212 552752 142218 552764
rect 143350 552752 143356 552764
rect 142212 552724 143356 552752
rect 142212 552712 142218 552724
rect 143350 552712 143356 552724
rect 143408 552712 143414 552764
rect 143534 552712 143540 552764
rect 143592 552752 143598 552764
rect 144730 552752 144736 552764
rect 143592 552724 144736 552752
rect 143592 552712 143598 552724
rect 144730 552712 144736 552724
rect 144788 552712 144794 552764
rect 144914 552712 144920 552764
rect 144972 552752 144978 552764
rect 146202 552752 146208 552764
rect 144972 552724 146208 552752
rect 144972 552712 144978 552724
rect 146202 552712 146208 552724
rect 146260 552712 146266 552764
rect 148502 552712 148508 552764
rect 148560 552752 148566 552764
rect 172514 552752 172520 552764
rect 148560 552724 172520 552752
rect 148560 552712 148566 552724
rect 172514 552712 172520 552724
rect 172572 552712 172578 552764
rect 179414 552712 179420 552764
rect 179472 552752 179478 552764
rect 180610 552752 180616 552764
rect 179472 552724 180616 552752
rect 179472 552712 179478 552724
rect 180610 552712 180616 552724
rect 180668 552712 180674 552764
rect 180886 552712 180892 552764
rect 180944 552752 180950 552764
rect 181990 552752 181996 552764
rect 180944 552724 181996 552752
rect 180944 552712 180950 552724
rect 181990 552712 181996 552724
rect 182048 552712 182054 552764
rect 190454 552712 190460 552764
rect 190512 552752 190518 552764
rect 191374 552752 191380 552764
rect 190512 552724 191380 552752
rect 190512 552712 190518 552724
rect 191374 552712 191380 552724
rect 191432 552712 191438 552764
rect 195974 552712 195980 552764
rect 196032 552752 196038 552764
rect 197078 552752 197084 552764
rect 196032 552724 197084 552752
rect 196032 552712 196038 552724
rect 197078 552712 197084 552724
rect 197136 552712 197142 552764
rect 198734 552712 198740 552764
rect 198792 552752 198798 552764
rect 199930 552752 199936 552764
rect 198792 552724 199936 552752
rect 198792 552712 198798 552724
rect 199930 552712 199936 552724
rect 199988 552712 199994 552764
rect 201494 552712 201500 552764
rect 201552 552752 201558 552764
rect 202782 552752 202788 552764
rect 201552 552724 202788 552752
rect 201552 552712 201558 552724
rect 202782 552712 202788 552724
rect 202840 552712 202846 552764
rect 213914 552712 213920 552764
rect 213972 552752 213978 552764
rect 215018 552752 215024 552764
rect 213972 552724 215024 552752
rect 213972 552712 213978 552724
rect 215018 552712 215024 552724
rect 215076 552712 215082 552764
rect 302510 552752 302516 552764
rect 215312 552724 302516 552752
rect 76800 552656 103652 552684
rect 76800 552644 76806 552656
rect 106274 552644 106280 552696
rect 106332 552684 106338 552696
rect 107562 552684 107568 552696
rect 106332 552656 107568 552684
rect 106332 552644 106338 552656
rect 107562 552644 107568 552656
rect 107620 552644 107626 552696
rect 110414 552644 110420 552696
rect 110472 552684 110478 552696
rect 111058 552684 111064 552696
rect 110472 552656 111064 552684
rect 110472 552644 110478 552656
rect 111058 552644 111064 552656
rect 111116 552644 111122 552696
rect 121822 552644 121828 552696
rect 121880 552644 121886 552696
rect 129734 552644 129740 552696
rect 129792 552644 129798 552696
rect 158714 552644 158720 552696
rect 158772 552684 158778 552696
rect 159818 552684 159824 552696
rect 158772 552656 159824 552684
rect 158772 552644 158778 552656
rect 159818 552644 159824 552656
rect 159876 552644 159882 552696
rect 212166 552644 212172 552696
rect 212224 552684 212230 552696
rect 215312 552684 215340 552724
rect 302510 552712 302516 552724
rect 302568 552712 302574 552764
rect 301314 552684 301320 552696
rect 212224 552656 215340 552684
rect 219406 552656 301320 552684
rect 212224 552644 212230 552656
rect 121454 552576 121460 552628
rect 121512 552616 121518 552628
rect 122558 552616 122564 552628
rect 121512 552588 122564 552616
rect 121512 552576 121518 552588
rect 122558 552576 122564 552588
rect 122616 552576 122622 552628
rect 210694 552576 210700 552628
rect 210752 552616 210758 552628
rect 219406 552616 219434 552656
rect 301314 552644 301320 552656
rect 301372 552644 301378 552696
rect 210752 552588 219434 552616
rect 210752 552576 210758 552588
rect 255314 552576 255320 552628
rect 255372 552616 255378 552628
rect 256510 552616 256516 552628
rect 255372 552588 256516 552616
rect 255372 552576 255378 552588
rect 256510 552576 256516 552588
rect 256568 552576 256574 552628
rect 266354 552576 266360 552628
rect 266412 552616 266418 552628
rect 267274 552616 267280 552628
rect 266412 552588 267280 552616
rect 266412 552576 266418 552588
rect 267274 552576 267280 552588
rect 267332 552576 267338 552628
rect 273254 552576 273260 552628
rect 273312 552616 273318 552628
rect 274450 552616 274456 552628
rect 273312 552588 274456 552616
rect 273312 552576 273318 552588
rect 274450 552576 274456 552588
rect 274508 552576 274514 552628
rect 293954 552576 293960 552628
rect 294012 552616 294018 552628
rect 295242 552616 295248 552628
rect 294012 552588 295248 552616
rect 294012 552576 294018 552588
rect 295242 552576 295248 552588
rect 295300 552576 295306 552628
rect 293126 552440 293132 552492
rect 293184 552480 293190 552492
rect 316954 552480 316960 552492
rect 293184 552452 316960 552480
rect 293184 552440 293190 552452
rect 316954 552440 316960 552452
rect 317012 552440 317018 552492
rect 290918 552372 290924 552424
rect 290976 552412 290982 552424
rect 316862 552412 316868 552424
rect 290976 552384 316868 552412
rect 290976 552372 290982 552384
rect 316862 552372 316868 552384
rect 316920 552372 316926 552424
rect 286686 552304 286692 552356
rect 286744 552344 286750 552356
rect 313918 552344 313924 552356
rect 286744 552316 313924 552344
rect 286744 552304 286750 552316
rect 313918 552304 313924 552316
rect 313976 552304 313982 552356
rect 285214 552236 285220 552288
rect 285272 552276 285278 552288
rect 317046 552276 317052 552288
rect 285272 552248 317052 552276
rect 285272 552236 285278 552248
rect 317046 552236 317052 552248
rect 317104 552236 317110 552288
rect 285950 552168 285956 552220
rect 286008 552208 286014 552220
rect 319438 552208 319444 552220
rect 286008 552180 319444 552208
rect 286008 552168 286014 552180
rect 319438 552168 319444 552180
rect 319496 552168 319502 552220
rect 252922 552100 252928 552152
rect 252980 552140 252986 552152
rect 322382 552140 322388 552152
rect 252980 552112 322388 552140
rect 252980 552100 252986 552112
rect 322382 552100 322388 552112
rect 322440 552100 322446 552152
rect 237926 552032 237932 552084
rect 237984 552072 237990 552084
rect 322566 552072 322572 552084
rect 237984 552044 322572 552072
rect 237984 552032 237990 552044
rect 322566 552032 322572 552044
rect 322624 552032 322630 552084
rect 148410 551964 148416 552016
rect 148468 552004 148474 552016
rect 149054 552004 149060 552016
rect 148468 551976 149060 552004
rect 148468 551964 148474 551976
rect 149054 551964 149060 551976
rect 149112 551964 149118 552016
rect 211430 551964 211436 552016
rect 211488 552004 211494 552016
rect 214650 552004 214656 552016
rect 211488 551976 214656 552004
rect 211488 551964 211494 551976
rect 214650 551964 214656 551976
rect 214708 551964 214714 552016
rect 148594 551896 148600 551948
rect 148652 551936 148658 551948
rect 149790 551936 149796 551948
rect 148652 551908 149796 551936
rect 148652 551896 148658 551908
rect 149790 551896 149796 551908
rect 149848 551896 149854 551948
rect 207106 551624 207112 551676
rect 207164 551664 207170 551676
rect 220262 551664 220268 551676
rect 207164 551636 220268 551664
rect 207164 551624 207170 551636
rect 220262 551624 220268 551636
rect 220320 551624 220326 551676
rect 207842 551556 207848 551608
rect 207900 551596 207906 551608
rect 229738 551596 229744 551608
rect 207900 551568 229744 551596
rect 207900 551556 207906 551568
rect 229738 551556 229744 551568
rect 229796 551556 229802 551608
rect 135438 551488 135444 551540
rect 135496 551528 135502 551540
rect 144270 551528 144276 551540
rect 135496 551500 144276 551528
rect 135496 551488 135502 551500
rect 144270 551488 144276 551500
rect 144328 551488 144334 551540
rect 147674 551488 147680 551540
rect 147732 551528 147738 551540
rect 191098 551528 191104 551540
rect 147732 551500 191104 551528
rect 147732 551488 147738 551500
rect 191098 551488 191104 551500
rect 191156 551488 191162 551540
rect 208578 551488 208584 551540
rect 208636 551528 208642 551540
rect 238294 551528 238300 551540
rect 208636 551500 238300 551528
rect 208636 551488 208642 551500
rect 238294 551488 238300 551500
rect 238352 551488 238358 551540
rect 152642 551420 152648 551472
rect 152700 551460 152706 551472
rect 211522 551460 211528 551472
rect 152700 551432 211528 551460
rect 152700 551420 152706 551432
rect 211522 551420 211528 551432
rect 211580 551420 211586 551472
rect 249426 551420 249432 551472
rect 249484 551460 249490 551472
rect 301498 551460 301504 551472
rect 249484 551432 301504 551460
rect 249484 551420 249490 551432
rect 301498 551420 301504 551432
rect 301556 551420 301562 551472
rect 120442 551352 120448 551404
rect 120500 551392 120506 551404
rect 130562 551392 130568 551404
rect 120500 551364 130568 551392
rect 120500 551352 120506 551364
rect 130562 551352 130568 551364
rect 130620 551352 130626 551404
rect 188522 551352 188528 551404
rect 188580 551392 188586 551404
rect 253934 551392 253940 551404
rect 188580 551364 253940 551392
rect 188580 551352 188586 551364
rect 253934 551352 253940 551364
rect 253992 551352 253998 551404
rect 57606 551284 57612 551336
rect 57664 551324 57670 551336
rect 77386 551324 77392 551336
rect 57664 551296 77392 551324
rect 57664 551284 57670 551296
rect 77386 551284 77392 551296
rect 77444 551284 77450 551336
rect 94590 551284 94596 551336
rect 94648 551324 94654 551336
rect 123386 551324 123392 551336
rect 94648 551296 123392 551324
rect 94648 551284 94654 551296
rect 123386 551284 123392 551296
rect 123444 551284 123450 551336
rect 124674 551284 124680 551336
rect 124732 551324 124738 551336
rect 210878 551324 210884 551336
rect 124732 551296 210884 551324
rect 124732 551284 124738 551296
rect 210878 551284 210884 551296
rect 210936 551284 210942 551336
rect 247218 551284 247224 551336
rect 247276 551324 247282 551336
rect 301590 551324 301596 551336
rect 247276 551296 301596 551324
rect 247276 551284 247282 551296
rect 301590 551284 301596 551296
rect 301648 551284 301654 551336
rect 265894 551216 265900 551268
rect 265952 551256 265958 551268
rect 307018 551256 307024 551268
rect 265952 551228 307024 551256
rect 265952 551216 265958 551228
rect 307018 551216 307024 551228
rect 307076 551216 307082 551268
rect 255866 551148 255872 551200
rect 255924 551188 255930 551200
rect 304442 551188 304448 551200
rect 255924 551160 304448 551188
rect 255924 551148 255930 551160
rect 304442 551148 304448 551160
rect 304500 551148 304506 551200
rect 273070 551080 273076 551132
rect 273128 551120 273134 551132
rect 321002 551120 321008 551132
rect 273128 551092 321008 551120
rect 273128 551080 273134 551092
rect 321002 551080 321008 551092
rect 321060 551080 321066 551132
rect 273714 551012 273720 551064
rect 273772 551052 273778 551064
rect 323762 551052 323768 551064
rect 273772 551024 323768 551052
rect 273772 551012 273778 551024
rect 323762 551012 323768 551024
rect 323820 551012 323826 551064
rect 265158 550944 265164 550996
rect 265216 550984 265222 550996
rect 318058 550984 318064 550996
rect 265216 550956 318064 550984
rect 265216 550944 265222 550956
rect 318058 550944 318064 550956
rect 318116 550944 318122 550996
rect 291654 550876 291660 550928
rect 291712 550916 291718 550928
rect 316770 550916 316776 550928
rect 291712 550888 316776 550916
rect 291712 550876 291718 550888
rect 316770 550876 316776 550888
rect 316828 550876 316834 550928
rect 287330 550808 287336 550860
rect 287388 550848 287394 550860
rect 317138 550848 317144 550860
rect 287388 550820 317144 550848
rect 287388 550808 287394 550820
rect 317138 550808 317144 550820
rect 317196 550808 317202 550860
rect 264422 550740 264428 550792
rect 264480 550780 264486 550792
rect 322474 550780 322480 550792
rect 264480 550752 322480 550780
rect 264480 550740 264486 550752
rect 322474 550740 322480 550752
rect 322532 550740 322538 550792
rect 263042 550672 263048 550724
rect 263100 550712 263106 550724
rect 322290 550712 322296 550724
rect 263100 550684 322296 550712
rect 263100 550672 263106 550684
rect 322290 550672 322296 550684
rect 322348 550672 322354 550724
rect 244366 550604 244372 550656
rect 244424 550644 244430 550656
rect 324866 550644 324872 550656
rect 244424 550616 324872 550644
rect 244424 550604 244430 550616
rect 324866 550604 324872 550616
rect 324924 550604 324930 550656
rect 84838 550536 84844 550588
rect 84896 550576 84902 550588
rect 86770 550576 86776 550588
rect 84896 550548 86776 550576
rect 84896 550536 84902 550548
rect 86770 550536 86776 550548
rect 86828 550536 86834 550588
rect 96062 550536 96068 550588
rect 96120 550576 96126 550588
rect 98638 550576 98644 550588
rect 96120 550548 98644 550576
rect 96120 550536 96126 550548
rect 98638 550536 98644 550548
rect 98696 550536 98702 550588
rect 104158 550536 104164 550588
rect 104216 550576 104222 550588
rect 105354 550576 105360 550588
rect 104216 550548 105360 550576
rect 104216 550536 104222 550548
rect 105354 550536 105360 550548
rect 105412 550536 105418 550588
rect 108298 550536 108304 550588
rect 108356 550576 108362 550588
rect 109678 550576 109684 550588
rect 108356 550548 109684 550576
rect 108356 550536 108362 550548
rect 109678 550536 109684 550548
rect 109736 550536 109742 550588
rect 115198 550536 115204 550588
rect 115256 550576 115262 550588
rect 116118 550576 116124 550588
rect 115256 550548 116124 550576
rect 115256 550536 115262 550548
rect 116118 550536 116124 550548
rect 116176 550536 116182 550588
rect 136174 550536 136180 550588
rect 136232 550576 136238 550588
rect 140038 550576 140044 550588
rect 136232 550548 140044 550576
rect 136232 550536 136238 550548
rect 140038 550536 140044 550548
rect 140096 550536 140102 550588
rect 146938 550536 146944 550588
rect 146996 550576 147002 550588
rect 148318 550576 148324 550588
rect 146996 550548 148324 550576
rect 146996 550536 147002 550548
rect 148318 550536 148324 550548
rect 148376 550536 148382 550588
rect 149882 550536 149888 550588
rect 149940 550576 149946 550588
rect 151262 550576 151268 550588
rect 149940 550548 151268 550576
rect 149940 550536 149946 550548
rect 151262 550536 151268 550548
rect 151320 550536 151326 550588
rect 230014 550536 230020 550588
rect 230072 550576 230078 550588
rect 231118 550576 231124 550588
rect 230072 550548 231124 550576
rect 230072 550536 230078 550548
rect 231118 550536 231124 550548
rect 231176 550536 231182 550588
rect 234338 550536 234344 550588
rect 234396 550576 234402 550588
rect 236638 550576 236644 550588
rect 234396 550548 236644 550576
rect 234396 550536 234402 550548
rect 236638 550536 236644 550548
rect 236696 550536 236702 550588
rect 291194 550536 291200 550588
rect 291252 550576 291258 550588
rect 292390 550576 292396 550588
rect 291252 550548 292396 550576
rect 291252 550536 291258 550548
rect 292390 550536 292396 550548
rect 292448 550536 292454 550588
rect 299566 550536 299572 550588
rect 299624 550576 299630 550588
rect 304350 550576 304356 550588
rect 299624 550548 304356 550576
rect 299624 550536 299630 550548
rect 304350 550536 304356 550548
rect 304408 550536 304414 550588
rect 55122 550468 55128 550520
rect 55180 550508 55186 550520
rect 67358 550508 67364 550520
rect 55180 550480 67364 550508
rect 55180 550468 55186 550480
rect 67358 550468 67364 550480
rect 67416 550468 67422 550520
rect 106918 550468 106924 550520
rect 106976 550508 106982 550520
rect 108942 550508 108948 550520
rect 106976 550480 108948 550508
rect 106976 550468 106982 550480
rect 108942 550468 108948 550480
rect 109000 550468 109006 550520
rect 298830 550468 298836 550520
rect 298888 550508 298894 550520
rect 304258 550508 304264 550520
rect 298888 550480 304264 550508
rect 298888 550468 298894 550480
rect 304258 550468 304264 550480
rect 304316 550468 304322 550520
rect 54938 550400 54944 550452
rect 54996 550440 55002 550452
rect 88886 550440 88892 550452
rect 54996 550412 88892 550440
rect 54996 550400 55002 550412
rect 88886 550400 88892 550412
rect 88944 550400 88950 550452
rect 91094 550400 91100 550452
rect 91152 550440 91158 550452
rect 96798 550440 96804 550452
rect 91152 550412 96804 550440
rect 91152 550400 91158 550412
rect 96798 550400 96804 550412
rect 96856 550400 96862 550452
rect 108390 550400 108396 550452
rect 108448 550440 108454 550452
rect 111794 550440 111800 550452
rect 108448 550412 111800 550440
rect 108448 550400 108454 550412
rect 111794 550400 111800 550412
rect 111852 550400 111858 550452
rect 171318 550400 171324 550452
rect 171376 550440 171382 550452
rect 173802 550440 173808 550452
rect 171376 550412 173808 550440
rect 171376 550400 171382 550412
rect 173802 550400 173808 550412
rect 173860 550400 173866 550452
rect 209222 550400 209228 550452
rect 209280 550440 209286 550452
rect 217318 550440 217324 550452
rect 209280 550412 217324 550440
rect 209280 550400 209286 550412
rect 217318 550400 217324 550412
rect 217376 550400 217382 550452
rect 58710 550332 58716 550384
rect 58768 550372 58774 550384
rect 95326 550372 95332 550384
rect 58768 550344 95332 550372
rect 58768 550332 58774 550344
rect 95326 550332 95332 550344
rect 95384 550332 95390 550384
rect 144086 550332 144092 550384
rect 144144 550372 144150 550384
rect 146294 550372 146300 550384
rect 144144 550344 146300 550372
rect 144144 550332 144150 550344
rect 146294 550332 146300 550344
rect 146352 550332 146358 550384
rect 151078 550332 151084 550384
rect 151136 550372 151142 550384
rect 153378 550372 153384 550384
rect 151136 550344 153384 550372
rect 151136 550332 151142 550344
rect 153378 550332 153384 550344
rect 153436 550332 153442 550384
rect 204254 550332 204260 550384
rect 204312 550372 204318 550384
rect 215938 550372 215944 550384
rect 204312 550344 215944 550372
rect 204312 550332 204318 550344
rect 215938 550332 215944 550344
rect 215996 550332 216002 550384
rect 56502 550264 56508 550316
rect 56560 550304 56566 550316
rect 83918 550304 83924 550316
rect 56560 550276 83924 550304
rect 56560 550264 56566 550276
rect 83918 550264 83924 550276
rect 83976 550264 83982 550316
rect 85298 550264 85304 550316
rect 85356 550304 85362 550316
rect 121638 550304 121644 550316
rect 85356 550276 121644 550304
rect 85356 550264 85362 550276
rect 121638 550264 121644 550276
rect 121696 550264 121702 550316
rect 157794 550264 157800 550316
rect 157852 550304 157858 550316
rect 166994 550304 167000 550316
rect 157852 550276 167000 550304
rect 157852 550264 157858 550276
rect 166994 550264 167000 550276
rect 167052 550264 167058 550316
rect 203518 550264 203524 550316
rect 203576 550304 203582 550316
rect 220078 550304 220084 550316
rect 203576 550276 220084 550304
rect 203576 550264 203582 550276
rect 220078 550264 220084 550276
rect 220136 550264 220142 550316
rect 225046 550264 225052 550316
rect 225104 550304 225110 550316
rect 235442 550304 235448 550316
rect 225104 550276 235448 550304
rect 225104 550264 225110 550276
rect 235442 550264 235448 550276
rect 235500 550264 235506 550316
rect 55030 550196 55036 550248
rect 55088 550236 55094 550248
rect 93210 550236 93216 550248
rect 55088 550208 93216 550236
rect 55088 550196 55094 550208
rect 93210 550196 93216 550208
rect 93268 550196 93274 550248
rect 114002 550196 114008 550248
rect 114060 550236 114066 550248
rect 125778 550236 125784 550248
rect 114060 550208 125784 550236
rect 114060 550196 114066 550208
rect 125778 550196 125784 550208
rect 125836 550196 125842 550248
rect 146110 550196 146116 550248
rect 146168 550236 146174 550248
rect 156966 550236 156972 550248
rect 146168 550208 156972 550236
rect 146168 550196 146174 550208
rect 156966 550196 156972 550208
rect 157024 550196 157030 550248
rect 169846 550196 169852 550248
rect 169904 550236 169910 550248
rect 175274 550236 175280 550248
rect 169904 550208 175280 550236
rect 169904 550196 169910 550208
rect 175274 550196 175280 550208
rect 175332 550196 175338 550248
rect 195606 550196 195612 550248
rect 195664 550236 195670 550248
rect 214558 550236 214564 550248
rect 195664 550208 214564 550236
rect 195664 550196 195670 550208
rect 214558 550196 214564 550208
rect 214616 550196 214622 550248
rect 219986 550196 219992 550248
rect 220044 550236 220050 550248
rect 233878 550236 233884 550248
rect 220044 550208 233884 550236
rect 220044 550196 220050 550208
rect 233878 550196 233884 550208
rect 233936 550196 233942 550248
rect 257246 550196 257252 550248
rect 257304 550236 257310 550248
rect 300578 550236 300584 550248
rect 257304 550208 300584 550236
rect 257304 550196 257310 550208
rect 300578 550196 300584 550208
rect 300636 550196 300642 550248
rect 56410 550128 56416 550180
rect 56468 550168 56474 550180
rect 98914 550168 98920 550180
rect 56468 550140 98920 550168
rect 56468 550128 56474 550140
rect 98914 550128 98920 550140
rect 98972 550128 98978 550180
rect 102778 550128 102784 550180
rect 102836 550168 102842 550180
rect 106090 550168 106096 550180
rect 102836 550140 106096 550168
rect 102836 550128 102842 550140
rect 106090 550128 106096 550140
rect 106148 550128 106154 550180
rect 106826 550128 106832 550180
rect 106884 550168 106890 550180
rect 124398 550168 124404 550180
rect 106884 550140 124404 550168
rect 106884 550128 106890 550140
rect 124398 550128 124404 550140
rect 124456 550128 124462 550180
rect 151998 550128 152004 550180
rect 152056 550168 152062 550180
rect 167730 550168 167736 550180
rect 152056 550140 167736 550168
rect 152056 550128 152062 550140
rect 167730 550128 167736 550140
rect 167788 550128 167794 550180
rect 170582 550128 170588 550180
rect 170640 550168 170646 550180
rect 195238 550168 195244 550180
rect 170640 550140 195244 550168
rect 170640 550128 170646 550140
rect 195238 550128 195244 550140
rect 195296 550128 195302 550180
rect 209958 550128 209964 550180
rect 210016 550168 210022 550180
rect 228358 550168 228364 550180
rect 210016 550140 228364 550168
rect 210016 550128 210022 550140
rect 228358 550128 228364 550140
rect 228416 550128 228422 550180
rect 230750 550128 230756 550180
rect 230808 550168 230814 550180
rect 244918 550168 244924 550180
rect 230808 550140 244924 550168
rect 230808 550128 230814 550140
rect 244918 550128 244924 550140
rect 244976 550128 244982 550180
rect 270862 550128 270868 550180
rect 270920 550168 270926 550180
rect 322750 550168 322756 550180
rect 270920 550140 322756 550168
rect 270920 550128 270926 550140
rect 322750 550128 322756 550140
rect 322808 550128 322814 550180
rect 57698 550060 57704 550112
rect 57756 550100 57762 550112
rect 99650 550100 99656 550112
rect 57756 550072 99656 550100
rect 57756 550060 57762 550072
rect 99650 550060 99656 550072
rect 99708 550060 99714 550112
rect 103974 550060 103980 550112
rect 104032 550100 104038 550112
rect 124306 550100 124312 550112
rect 104032 550072 124312 550100
rect 104032 550060 104038 550072
rect 124306 550060 124312 550072
rect 124364 550060 124370 550112
rect 139026 550060 139032 550112
rect 139084 550100 139090 550112
rect 184290 550100 184296 550112
rect 139084 550072 184296 550100
rect 139084 550060 139090 550072
rect 184290 550060 184296 550072
rect 184348 550060 184354 550112
rect 194226 550060 194232 550112
rect 194284 550100 194290 550112
rect 220170 550100 220176 550112
rect 194284 550072 220176 550100
rect 194284 550060 194290 550072
rect 220170 550060 220176 550072
rect 220228 550060 220234 550112
rect 225782 550060 225788 550112
rect 225840 550100 225846 550112
rect 241514 550100 241520 550112
rect 225840 550072 241520 550100
rect 225840 550060 225846 550072
rect 241514 550060 241520 550072
rect 241572 550060 241578 550112
rect 242250 550060 242256 550112
rect 242308 550100 242314 550112
rect 323946 550100 323952 550112
rect 242308 550072 323952 550100
rect 242308 550060 242314 550072
rect 323946 550060 323952 550072
rect 324004 550060 324010 550112
rect 56318 549992 56324 550044
rect 56376 550032 56382 550044
rect 73798 550032 73804 550044
rect 56376 550004 73804 550032
rect 56376 549992 56382 550004
rect 73798 549992 73804 550004
rect 73856 549992 73862 550044
rect 78122 549992 78128 550044
rect 78180 550032 78186 550044
rect 122190 550032 122196 550044
rect 78180 550004 122196 550032
rect 78180 549992 78186 550004
rect 122190 549992 122196 550004
rect 122248 549992 122254 550044
rect 136910 549992 136916 550044
rect 136968 550032 136974 550044
rect 156598 550032 156604 550044
rect 136968 550004 156604 550032
rect 136968 549992 136974 550004
rect 156598 549992 156604 550004
rect 156656 549992 156662 550044
rect 160094 549992 160100 550044
rect 160152 550032 160158 550044
rect 172698 550032 172704 550044
rect 160152 550004 172704 550032
rect 160152 549992 160158 550004
rect 172698 549992 172704 550004
rect 172756 549992 172762 550044
rect 183462 549992 183468 550044
rect 183520 550032 183526 550044
rect 231210 550032 231216 550044
rect 183520 550004 231216 550032
rect 183520 549992 183526 550004
rect 231210 549992 231216 550004
rect 231268 549992 231274 550044
rect 60366 549924 60372 549976
rect 60424 549964 60430 549976
rect 116854 549964 116860 549976
rect 60424 549936 116860 549964
rect 60424 549924 60430 549936
rect 116854 549924 116860 549936
rect 116912 549924 116918 549976
rect 128998 549924 129004 549976
rect 129056 549964 129062 549976
rect 137186 549964 137192 549976
rect 129056 549936 137192 549964
rect 129056 549924 129062 549936
rect 137186 549924 137192 549936
rect 137244 549924 137250 549976
rect 154114 549924 154120 549976
rect 154172 549964 154178 549976
rect 204898 549964 204904 549976
rect 154172 549936 204904 549964
rect 154172 549924 154178 549936
rect 204898 549924 204904 549936
rect 204956 549924 204962 549976
rect 212810 549924 212816 549976
rect 212868 549964 212874 549976
rect 249058 549964 249064 549976
rect 212868 549936 249064 549964
rect 212868 549924 212874 549936
rect 249058 549924 249064 549936
rect 249116 549924 249122 549976
rect 252278 549924 252284 549976
rect 252336 549964 252342 549976
rect 293954 549964 293960 549976
rect 252336 549936 293960 549964
rect 252336 549924 252342 549936
rect 293954 549924 293960 549936
rect 294012 549924 294018 549976
rect 58618 549856 58624 549908
rect 58676 549896 58682 549908
rect 117590 549896 117596 549908
rect 58676 549868 117596 549896
rect 58676 549856 58682 549868
rect 117590 549856 117596 549868
rect 117648 549856 117654 549908
rect 118970 549856 118976 549908
rect 119028 549896 119034 549908
rect 128906 549896 128912 549908
rect 119028 549868 128912 549896
rect 119028 549856 119034 549868
rect 128906 549856 128912 549868
rect 128964 549856 128970 549908
rect 131850 549856 131856 549908
rect 131908 549896 131914 549908
rect 144178 549896 144184 549908
rect 131908 549868 144184 549896
rect 131908 549856 131914 549868
rect 144178 549856 144184 549868
rect 144236 549856 144242 549908
rect 148962 549856 148968 549908
rect 149020 549896 149026 549908
rect 171962 549896 171968 549908
rect 149020 549868 171968 549896
rect 149020 549856 149026 549868
rect 171962 549856 171968 549868
rect 172020 549856 172026 549908
rect 176286 549856 176292 549908
rect 176344 549896 176350 549908
rect 238110 549896 238116 549908
rect 176344 549868 238116 549896
rect 176344 549856 176350 549868
rect 238110 549856 238116 549868
rect 238168 549856 238174 549908
rect 280154 549856 280160 549908
rect 280212 549896 280218 549908
rect 301682 549896 301688 549908
rect 280212 549868 301688 549896
rect 280212 549856 280218 549868
rect 301682 549856 301688 549868
rect 301740 549856 301746 549908
rect 169754 549788 169760 549840
rect 169812 549828 169818 549840
rect 173434 549828 173440 549840
rect 169812 549800 173440 549828
rect 169812 549788 169818 549800
rect 173434 549788 173440 549800
rect 173492 549788 173498 549840
rect 276566 549788 276572 549840
rect 276624 549828 276630 549840
rect 300118 549828 300124 549840
rect 276624 549800 300124 549828
rect 276624 549788 276630 549800
rect 300118 549788 300124 549800
rect 300176 549788 300182 549840
rect 277302 549720 277308 549772
rect 277360 549760 277366 549772
rect 300394 549760 300400 549772
rect 277360 549732 300400 549760
rect 277360 549720 277366 549732
rect 300394 549720 300400 549732
rect 300452 549720 300458 549772
rect 275922 549652 275928 549704
rect 275980 549692 275986 549704
rect 302878 549692 302884 549704
rect 275980 549664 302884 549692
rect 275980 549652 275986 549664
rect 302878 549652 302884 549664
rect 302936 549652 302942 549704
rect 284478 549584 284484 549636
rect 284536 549624 284542 549636
rect 319530 549624 319536 549636
rect 284536 549596 319536 549624
rect 284536 549584 284542 549596
rect 319530 549584 319536 549596
rect 319588 549584 319594 549636
rect 294506 549516 294512 549568
rect 294564 549556 294570 549568
rect 319714 549556 319720 549568
rect 294564 549528 319720 549556
rect 294564 549516 294570 549528
rect 319714 549516 319720 549528
rect 319772 549516 319778 549568
rect 243630 549448 243636 549500
rect 243688 549488 243694 549500
rect 287606 549488 287612 549500
rect 243688 549460 287612 549488
rect 243688 549448 243694 549460
rect 287606 549448 287612 549460
rect 287664 549448 287670 549500
rect 289786 549460 292574 549488
rect 109770 549380 109776 549432
rect 109828 549420 109834 549432
rect 114646 549420 114652 549432
rect 109828 549392 114652 549420
rect 109828 549380 109834 549392
rect 114646 549380 114652 549392
rect 114704 549380 114710 549432
rect 283098 549380 283104 549432
rect 283156 549420 283162 549432
rect 289786 549420 289814 549460
rect 283156 549392 289814 549420
rect 292546 549420 292574 549460
rect 295978 549448 295984 549500
rect 296036 549488 296042 549500
rect 319622 549488 319628 549500
rect 296036 549460 319628 549488
rect 296036 549448 296042 549460
rect 319622 549448 319628 549460
rect 319680 549448 319686 549500
rect 322658 549420 322664 549432
rect 292546 549392 322664 549420
rect 283156 549380 283162 549392
rect 322658 549380 322664 549392
rect 322716 549380 322722 549432
rect 61654 549312 61660 549364
rect 61712 549352 61718 549364
rect 64966 549352 64972 549364
rect 61712 549324 64972 549352
rect 61712 549312 61718 549324
rect 64966 549312 64972 549324
rect 65024 549312 65030 549364
rect 118234 549312 118240 549364
rect 118292 549352 118298 549364
rect 124858 549352 124864 549364
rect 118292 549324 124864 549352
rect 118292 549312 118298 549324
rect 124858 549312 124864 549324
rect 124916 549312 124922 549364
rect 287882 549312 287888 549364
rect 287940 549352 287946 549364
rect 300486 549352 300492 549364
rect 287940 549324 300492 549352
rect 287940 549312 287946 549324
rect 300486 549312 300492 549324
rect 300544 549312 300550 549364
rect 278038 549244 278044 549296
rect 278096 549284 278102 549296
rect 300302 549284 300308 549296
rect 278096 549256 300308 549284
rect 278096 549244 278102 549256
rect 300302 549244 300308 549256
rect 300360 549244 300366 549296
rect 296714 548768 296720 548820
rect 296772 548808 296778 548820
rect 319806 548808 319812 548820
rect 296772 548780 319812 548808
rect 296772 548768 296778 548780
rect 319806 548768 319812 548780
rect 319864 548768 319870 548820
rect 278774 548700 278780 548752
rect 278832 548740 278838 548752
rect 300762 548740 300768 548752
rect 278832 548712 300768 548740
rect 278832 548700 278838 548712
rect 300762 548700 300768 548712
rect 300820 548700 300826 548752
rect 281626 548632 281632 548684
rect 281684 548672 281690 548684
rect 287882 548672 287888 548684
rect 281684 548644 287888 548672
rect 281684 548632 281690 548644
rect 287882 548632 287888 548644
rect 287940 548632 287946 548684
rect 293954 548632 293960 548684
rect 294012 548672 294018 548684
rect 321830 548672 321836 548684
rect 294012 548644 321836 548672
rect 294012 548632 294018 548644
rect 321830 548632 321836 548644
rect 321888 548632 321894 548684
rect 268746 548564 268752 548616
rect 268804 548604 268810 548616
rect 300210 548604 300216 548616
rect 268804 548576 300216 548604
rect 268804 548564 268810 548576
rect 300210 548564 300216 548576
rect 300268 548564 300274 548616
rect 287606 548496 287612 548548
rect 287664 548536 287670 548548
rect 322198 548536 322204 548548
rect 287664 548508 322204 548536
rect 287664 548496 287670 548508
rect 322198 548496 322204 548508
rect 322256 548496 322262 548548
rect 272334 548428 272340 548480
rect 272392 548468 272398 548480
rect 304258 548468 304264 548480
rect 272392 548440 304264 548468
rect 272392 548428 272398 548440
rect 304258 548428 304264 548440
rect 304316 548428 304322 548480
rect 262306 548360 262312 548412
rect 262364 548400 262370 548412
rect 324774 548400 324780 548412
rect 262364 548372 324780 548400
rect 262364 548360 262370 548372
rect 324774 548360 324780 548372
rect 324832 548360 324838 548412
rect 260834 548292 260840 548344
rect 260892 548332 260898 548344
rect 323670 548332 323676 548344
rect 260892 548304 323676 548332
rect 260892 548292 260898 548304
rect 323670 548292 323676 548304
rect 323728 548292 323734 548344
rect 240042 548224 240048 548276
rect 240100 548264 240106 548276
rect 302970 548264 302976 548276
rect 240100 548236 302976 548264
rect 240100 548224 240106 548236
rect 302970 548224 302976 548236
rect 303028 548224 303034 548276
rect 236454 548156 236460 548208
rect 236512 548196 236518 548208
rect 302050 548196 302056 548208
rect 236512 548168 302056 548196
rect 236512 548156 236518 548168
rect 302050 548156 302056 548168
rect 302108 548156 302114 548208
rect 235810 548088 235816 548140
rect 235868 548088 235874 548140
rect 254394 548088 254400 548140
rect 254452 548128 254458 548140
rect 324682 548128 324688 548140
rect 254452 548100 324688 548128
rect 254452 548088 254458 548100
rect 324682 548088 324688 548100
rect 324740 548088 324746 548140
rect 235828 548060 235856 548088
rect 323854 548060 323860 548072
rect 235828 548032 323860 548060
rect 323854 548020 323860 548032
rect 323912 548020 323918 548072
rect 300762 542308 300768 542360
rect 300820 542348 300826 542360
rect 321554 542348 321560 542360
rect 300820 542320 321560 542348
rect 300820 542308 300826 542320
rect 321554 542308 321560 542320
rect 321612 542308 321618 542360
rect 302602 539588 302608 539640
rect 302660 539628 302666 539640
rect 320818 539628 320824 539640
rect 302660 539600 320824 539628
rect 302660 539588 302666 539600
rect 320818 539588 320824 539600
rect 320876 539588 320882 539640
rect 302050 536732 302056 536784
rect 302108 536772 302114 536784
rect 321554 536772 321560 536784
rect 302108 536744 321560 536772
rect 302108 536732 302114 536744
rect 321554 536732 321560 536744
rect 321612 536732 321618 536784
rect 436738 527960 436744 528012
rect 436796 528000 436802 528012
rect 436922 528000 436928 528012
rect 436796 527972 436928 528000
rect 436796 527960 436802 527972
rect 436922 527960 436928 527972
rect 436980 527960 436986 528012
rect 436370 527688 436376 527740
rect 436428 527728 436434 527740
rect 436646 527728 436652 527740
rect 436428 527700 436652 527728
rect 436428 527688 436434 527700
rect 436646 527688 436652 527700
rect 436704 527688 436710 527740
rect 302970 527076 302976 527128
rect 303028 527116 303034 527128
rect 321554 527116 321560 527128
rect 303028 527088 321560 527116
rect 303028 527076 303034 527088
rect 321554 527076 321560 527088
rect 321612 527076 321618 527128
rect 300486 522928 300492 522980
rect 300544 522968 300550 522980
rect 436554 522968 436560 522980
rect 300544 522940 436560 522968
rect 300544 522928 300550 522940
rect 436554 522928 436560 522940
rect 436612 522928 436618 522980
rect 300394 522860 300400 522912
rect 300452 522900 300458 522912
rect 436462 522900 436468 522912
rect 300452 522872 436468 522900
rect 300452 522860 300458 522872
rect 436462 522860 436468 522872
rect 436520 522860 436526 522912
rect 300578 522792 300584 522844
rect 300636 522832 300642 522844
rect 436186 522832 436192 522844
rect 300636 522804 436192 522832
rect 300636 522792 300642 522804
rect 436186 522792 436192 522804
rect 436244 522792 436250 522844
rect 301774 522724 301780 522776
rect 301832 522764 301838 522776
rect 436830 522764 436836 522776
rect 301832 522736 436836 522764
rect 301832 522724 301838 522736
rect 436830 522724 436836 522736
rect 436888 522724 436894 522776
rect 301866 522656 301872 522708
rect 301924 522696 301930 522708
rect 433518 522696 433524 522708
rect 301924 522668 433524 522696
rect 301924 522656 301930 522668
rect 433518 522656 433524 522668
rect 433576 522656 433582 522708
rect 321094 522588 321100 522640
rect 321152 522628 321158 522640
rect 436094 522628 436100 522640
rect 321152 522600 436100 522628
rect 321152 522588 321158 522600
rect 436094 522588 436100 522600
rect 436152 522588 436158 522640
rect 322750 522520 322756 522572
rect 322808 522560 322814 522572
rect 436646 522560 436652 522572
rect 322808 522532 436652 522560
rect 322808 522520 322814 522532
rect 436646 522520 436652 522532
rect 436704 522520 436710 522572
rect 323946 522452 323952 522504
rect 324004 522492 324010 522504
rect 436738 522492 436744 522504
rect 324004 522464 436744 522492
rect 324004 522452 324010 522464
rect 436738 522452 436744 522464
rect 436796 522452 436802 522504
rect 324866 522384 324872 522436
rect 324924 522424 324930 522436
rect 325142 522424 325148 522436
rect 324924 522396 325148 522424
rect 324924 522384 324930 522396
rect 325142 522384 325148 522396
rect 325200 522384 325206 522436
rect 323578 521568 323584 521620
rect 323636 521608 323642 521620
rect 342714 521608 342720 521620
rect 323636 521580 342720 521608
rect 323636 521568 323642 521580
rect 342714 521568 342720 521580
rect 342772 521568 342778 521620
rect 319438 521500 319444 521552
rect 319496 521540 319502 521552
rect 495434 521540 495440 521552
rect 319496 521512 495440 521540
rect 319496 521500 319502 521512
rect 495434 521500 495440 521512
rect 495492 521500 495498 521552
rect 319806 521432 319812 521484
rect 319864 521472 319870 521484
rect 459554 521472 459560 521484
rect 319864 521444 459560 521472
rect 319864 521432 319870 521444
rect 459554 521432 459560 521444
rect 459612 521432 459618 521484
rect 319622 521364 319628 521416
rect 319680 521404 319686 521416
rect 457438 521404 457444 521416
rect 319680 521376 457444 521404
rect 319680 521364 319686 521376
rect 457438 521364 457444 521376
rect 457496 521364 457502 521416
rect 300302 521296 300308 521348
rect 300360 521336 300366 521348
rect 436922 521336 436928 521348
rect 300360 521308 436928 521336
rect 300360 521296 300366 521308
rect 436922 521296 436928 521308
rect 436980 521296 436986 521348
rect 301682 521228 301688 521280
rect 301740 521268 301746 521280
rect 436278 521268 436284 521280
rect 301740 521240 436284 521268
rect 301740 521228 301746 521240
rect 436278 521228 436284 521240
rect 436336 521228 436342 521280
rect 300118 521160 300124 521212
rect 300176 521200 300182 521212
rect 419994 521200 420000 521212
rect 300176 521172 420000 521200
rect 300176 521160 300182 521172
rect 419994 521160 420000 521172
rect 420052 521160 420058 521212
rect 319530 521092 319536 521144
rect 319588 521132 319594 521144
rect 433426 521132 433432 521144
rect 319588 521104 433432 521132
rect 319588 521092 319594 521104
rect 433426 521092 433432 521104
rect 433484 521092 433490 521144
rect 322382 521024 322388 521076
rect 322440 521064 322446 521076
rect 433702 521064 433708 521076
rect 322440 521036 433708 521064
rect 322440 521024 322446 521036
rect 433702 521024 433708 521036
rect 433760 521024 433766 521076
rect 322566 520956 322572 521008
rect 322624 520996 322630 521008
rect 433610 520996 433616 521008
rect 322624 520968 433616 520996
rect 322624 520956 322630 520968
rect 433610 520956 433616 520968
rect 433668 520956 433674 521008
rect 322658 520888 322664 520940
rect 322716 520928 322722 520940
rect 433334 520928 433340 520940
rect 322716 520900 433340 520928
rect 322716 520888 322722 520900
rect 433334 520888 433340 520900
rect 433392 520888 433398 520940
rect 305638 520820 305644 520872
rect 305696 520860 305702 520872
rect 374270 520860 374276 520872
rect 305696 520832 374276 520860
rect 305696 520820 305702 520832
rect 374270 520820 374276 520832
rect 374328 520820 374334 520872
rect 302878 520752 302884 520804
rect 302936 520792 302942 520804
rect 356238 520792 356244 520804
rect 302936 520764 356244 520792
rect 302936 520752 302942 520764
rect 356238 520752 356244 520764
rect 356296 520752 356302 520804
rect 319714 520684 319720 520736
rect 319772 520724 319778 520736
rect 500954 520724 500960 520736
rect 319772 520696 500960 520724
rect 319772 520684 319778 520696
rect 500954 520684 500960 520696
rect 501012 520684 501018 520736
rect 323670 520276 323676 520328
rect 323728 520316 323734 520328
rect 323728 520288 324820 520316
rect 323728 520276 323734 520288
rect 318058 520208 318064 520260
rect 318116 520248 318122 520260
rect 324682 520248 324688 520260
rect 318116 520220 324688 520248
rect 318116 520208 318122 520220
rect 324682 520208 324688 520220
rect 324740 520208 324746 520260
rect 324792 520248 324820 520288
rect 347222 520248 347228 520260
rect 324792 520220 347228 520248
rect 347222 520208 347228 520220
rect 347280 520208 347286 520260
rect 323854 520140 323860 520192
rect 323912 520180 323918 520192
rect 338206 520180 338212 520192
rect 323912 520152 338212 520180
rect 323912 520140 323918 520152
rect 338206 520140 338212 520152
rect 338264 520140 338270 520192
rect 324590 520072 324596 520124
rect 324648 520112 324654 520124
rect 334066 520112 334072 520124
rect 324648 520084 334072 520112
rect 324648 520072 324654 520084
rect 334066 520072 334072 520084
rect 334124 520072 334130 520124
rect 300210 520004 300216 520056
rect 300268 520044 300274 520056
rect 393314 520044 393320 520056
rect 300268 520016 393320 520044
rect 300268 520004 300274 520016
rect 393314 520004 393320 520016
rect 393372 520004 393378 520056
rect 322290 519936 322296 519988
rect 322348 519976 322354 519988
rect 406470 519976 406476 519988
rect 322348 519948 406476 519976
rect 322348 519936 322354 519948
rect 406470 519936 406476 519948
rect 406528 519936 406534 519988
rect 307018 519868 307024 519920
rect 307076 519908 307082 519920
rect 388438 519908 388444 519920
rect 307076 519880 388444 519908
rect 307076 519868 307082 519880
rect 388438 519868 388444 519880
rect 388496 519868 388502 519920
rect 323762 519800 323768 519852
rect 323820 519840 323826 519852
rect 401962 519840 401968 519852
rect 323820 519812 401968 519840
rect 323820 519800 323826 519812
rect 401962 519800 401968 519812
rect 402020 519800 402026 519852
rect 301590 519732 301596 519784
rect 301648 519772 301654 519784
rect 365254 519772 365260 519784
rect 301648 519744 365260 519772
rect 301648 519732 301654 519744
rect 365254 519732 365260 519744
rect 365312 519732 365318 519784
rect 322474 519664 322480 519716
rect 322532 519704 322538 519716
rect 379514 519704 379520 519716
rect 322532 519676 379520 519704
rect 322532 519664 322538 519676
rect 379514 519664 379520 519676
rect 379572 519664 379578 519716
rect 321002 519596 321008 519648
rect 321060 519636 321066 519648
rect 369854 519636 369860 519648
rect 321060 519608 369860 519636
rect 321060 519596 321066 519608
rect 369854 519596 369860 519608
rect 369912 519596 369918 519648
rect 324498 519528 324504 519580
rect 324556 519568 324562 519580
rect 351914 519568 351920 519580
rect 324556 519540 351920 519568
rect 324556 519528 324562 519540
rect 351914 519528 351920 519540
rect 351972 519528 351978 519580
rect 304258 519460 304264 519512
rect 304316 519500 304322 519512
rect 415486 519500 415492 519512
rect 304316 519472 415492 519500
rect 304316 519460 304322 519472
rect 415486 519460 415492 519472
rect 415544 519460 415550 519512
rect 304442 519392 304448 519444
rect 304500 519432 304506 519444
rect 411346 519432 411352 519444
rect 304500 519404 411352 519432
rect 304500 519392 304506 519404
rect 411346 519392 411352 519404
rect 411404 519392 411410 519444
rect 325142 519324 325148 519376
rect 325200 519364 325206 519376
rect 424502 519364 424508 519376
rect 325200 519336 424508 519364
rect 325200 519324 325206 519336
rect 424502 519324 424508 519336
rect 424560 519324 424566 519376
rect 317138 518848 317144 518900
rect 317196 518888 317202 518900
rect 476114 518888 476120 518900
rect 317196 518860 476120 518888
rect 317196 518848 317202 518860
rect 476114 518848 476120 518860
rect 476172 518848 476178 518900
rect 317046 518780 317052 518832
rect 317104 518820 317110 518832
rect 470594 518820 470600 518832
rect 317104 518792 470600 518820
rect 317104 518780 317110 518792
rect 470594 518780 470600 518792
rect 470652 518780 470658 518832
rect 316770 518712 316776 518764
rect 316828 518752 316834 518764
rect 457622 518752 457628 518764
rect 316828 518724 457628 518752
rect 316828 518712 316834 518724
rect 457622 518712 457628 518724
rect 457680 518712 457686 518764
rect 302970 518168 302976 518220
rect 303028 518208 303034 518220
rect 576118 518208 576124 518220
rect 303028 518180 576124 518208
rect 303028 518168 303034 518180
rect 576118 518168 576124 518180
rect 576176 518168 576182 518220
rect 52362 517488 52368 517540
rect 52420 517528 52426 517540
rect 57882 517528 57888 517540
rect 52420 517500 57888 517528
rect 52420 517488 52426 517500
rect 57882 517488 57888 517500
rect 57940 517488 57946 517540
rect 313918 517420 313924 517472
rect 313976 517460 313982 517472
rect 512178 517460 512184 517472
rect 313976 517432 512184 517460
rect 313976 517420 313982 517432
rect 512178 517420 512184 517432
rect 512236 517420 512242 517472
rect 316954 517352 316960 517404
rect 317012 517392 317018 517404
rect 512270 517392 512276 517404
rect 317012 517364 512276 517392
rect 317012 517352 317018 517364
rect 512270 517352 512276 517364
rect 512328 517352 512334 517404
rect 316862 517284 316868 517336
rect 316920 517324 316926 517336
rect 488534 517324 488540 517336
rect 316920 517296 488540 517324
rect 316920 517284 316926 517296
rect 488534 517284 488540 517296
rect 488592 517284 488598 517336
rect 317230 517216 317236 517268
rect 317288 517256 317294 517268
rect 465074 517256 465080 517268
rect 317288 517228 465080 517256
rect 317288 517216 317294 517228
rect 465074 517216 465080 517228
rect 465132 517216 465138 517268
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 11698 514808 11704 514820
rect 3476 514780 11704 514808
rect 3476 514768 3482 514780
rect 11698 514768 11704 514780
rect 11756 514768 11762 514820
rect 560938 511912 560944 511964
rect 560996 511952 561002 511964
rect 580166 511952 580172 511964
rect 560996 511924 580172 511952
rect 560996 511912 561002 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 302234 495456 302240 495508
rect 302292 495496 302298 495508
rect 520918 495496 520924 495508
rect 302292 495468 520924 495496
rect 302292 495456 302298 495468
rect 520918 495456 520924 495468
rect 520976 495456 520982 495508
rect 320818 489132 320824 489184
rect 320876 489172 320882 489184
rect 580258 489172 580264 489184
rect 320876 489144 580264 489172
rect 320876 489132 320882 489144
rect 580258 489132 580264 489144
rect 580316 489132 580322 489184
rect 11698 488044 11704 488096
rect 11756 488084 11762 488096
rect 360194 488084 360200 488096
rect 11756 488056 360200 488084
rect 11756 488044 11762 488056
rect 360194 488044 360200 488056
rect 360252 488044 360258 488096
rect 293970 487772 293976 487824
rect 294028 487812 294034 487824
rect 294138 487812 294144 487824
rect 294028 487784 294144 487812
rect 294028 487772 294034 487784
rect 294138 487772 294144 487784
rect 294196 487772 294202 487824
rect 205818 487024 205824 487076
rect 205876 487064 205882 487076
rect 206094 487064 206100 487076
rect 205876 487036 206100 487064
rect 205876 487024 205882 487036
rect 206094 487024 206100 487036
rect 206152 487024 206158 487076
rect 109494 486616 109500 486668
rect 109552 486656 109558 486668
rect 204254 486656 204260 486668
rect 109552 486628 204260 486656
rect 109552 486616 109558 486628
rect 204254 486616 204260 486628
rect 204312 486616 204318 486668
rect 109402 486548 109408 486600
rect 109460 486588 109466 486600
rect 205634 486588 205640 486600
rect 109460 486560 205640 486588
rect 109460 486548 109466 486560
rect 205634 486548 205640 486560
rect 205692 486548 205698 486600
rect 51902 486480 51908 486532
rect 51960 486520 51966 486532
rect 99374 486520 99380 486532
rect 51960 486492 99380 486520
rect 51960 486480 51966 486492
rect 99374 486480 99380 486492
rect 99432 486480 99438 486532
rect 140866 486480 140872 486532
rect 140924 486520 140930 486532
rect 199102 486520 199108 486532
rect 140924 486492 199108 486520
rect 140924 486480 140930 486492
rect 199102 486480 199108 486492
rect 199160 486480 199166 486532
rect 203610 486480 203616 486532
rect 203668 486520 203674 486532
rect 356606 486520 356612 486532
rect 203668 486492 356612 486520
rect 203668 486480 203674 486492
rect 356606 486480 356612 486492
rect 356664 486480 356670 486532
rect 15838 486412 15844 486464
rect 15896 486452 15902 486464
rect 383654 486452 383660 486464
rect 15896 486424 383660 486452
rect 15896 486412 15902 486424
rect 383654 486412 383660 486424
rect 383712 486412 383718 486464
rect 56410 485732 56416 485784
rect 56468 485772 56474 485784
rect 81710 485772 81716 485784
rect 56468 485744 81716 485772
rect 56468 485732 56474 485744
rect 81710 485732 81716 485744
rect 81768 485732 81774 485784
rect 151262 485732 151268 485784
rect 151320 485772 151326 485784
rect 211154 485772 211160 485784
rect 151320 485744 211160 485772
rect 151320 485732 151326 485744
rect 211154 485732 211160 485744
rect 211212 485732 211218 485784
rect 73890 485664 73896 485716
rect 73948 485704 73954 485716
rect 102870 485704 102876 485716
rect 73948 485676 102876 485704
rect 73948 485664 73954 485676
rect 102870 485664 102876 485676
rect 102928 485664 102934 485716
rect 153930 485664 153936 485716
rect 153988 485704 153994 485716
rect 212534 485704 212540 485716
rect 153988 485676 212540 485704
rect 153988 485664 153994 485676
rect 212534 485664 212540 485676
rect 212592 485664 212598 485716
rect 59906 485596 59912 485648
rect 59964 485636 59970 485648
rect 91830 485636 91836 485648
rect 59964 485608 91836 485636
rect 59964 485596 59970 485608
rect 91830 485596 91836 485608
rect 91888 485596 91894 485648
rect 166166 485596 166172 485648
rect 166224 485636 166230 485648
rect 211154 485636 211160 485648
rect 166224 485608 211160 485636
rect 166224 485596 166230 485608
rect 211154 485596 211160 485608
rect 211212 485596 211218 485648
rect 56502 485528 56508 485580
rect 56560 485568 56566 485580
rect 89162 485568 89168 485580
rect 56560 485540 89168 485568
rect 56560 485528 56566 485540
rect 89162 485528 89168 485540
rect 89220 485528 89226 485580
rect 150434 485528 150440 485580
rect 150492 485568 150498 485580
rect 150492 485540 201356 485568
rect 150492 485528 150498 485540
rect 69658 485460 69664 485512
rect 69716 485500 69722 485512
rect 92290 485500 92296 485512
rect 69716 485472 92296 485500
rect 69716 485460 69722 485472
rect 92290 485460 92296 485472
rect 92348 485460 92354 485512
rect 152182 485460 152188 485512
rect 152240 485500 152246 485512
rect 201328 485500 201356 485540
rect 201402 485528 201408 485580
rect 201460 485568 201466 485580
rect 211614 485568 211620 485580
rect 201460 485540 211620 485568
rect 201460 485528 201466 485540
rect 211614 485528 211620 485540
rect 211672 485528 211678 485580
rect 242066 485528 242072 485580
rect 242124 485568 242130 485580
rect 356698 485568 356704 485580
rect 242124 485540 356704 485568
rect 242124 485528 242130 485540
rect 356698 485528 356704 485540
rect 356756 485528 356762 485580
rect 206186 485500 206192 485512
rect 152240 485472 201264 485500
rect 201328 485472 206192 485500
rect 152240 485460 152246 485472
rect 56318 485392 56324 485444
rect 56376 485432 56382 485444
rect 88334 485432 88340 485444
rect 56376 485404 88340 485432
rect 56376 485392 56382 485404
rect 88334 485392 88340 485404
rect 88392 485392 88398 485444
rect 149422 485392 149428 485444
rect 149480 485432 149486 485444
rect 191190 485432 191196 485444
rect 149480 485404 191196 485432
rect 149480 485392 149486 485404
rect 191190 485392 191196 485404
rect 191248 485392 191254 485444
rect 201236 485432 201264 485472
rect 206186 485460 206192 485472
rect 206244 485460 206250 485512
rect 240042 485460 240048 485512
rect 240100 485500 240106 485512
rect 358262 485500 358268 485512
rect 240100 485472 358268 485500
rect 240100 485460 240106 485472
rect 358262 485460 358268 485472
rect 358320 485460 358326 485512
rect 204438 485432 204444 485444
rect 201236 485404 204444 485432
rect 204438 485392 204444 485404
rect 204496 485392 204502 485444
rect 208302 485392 208308 485444
rect 208360 485432 208366 485444
rect 217410 485432 217416 485444
rect 208360 485404 217416 485432
rect 208360 485392 208366 485404
rect 217410 485392 217416 485404
rect 217468 485392 217474 485444
rect 239674 485392 239680 485444
rect 239732 485432 239738 485444
rect 358354 485432 358360 485444
rect 239732 485404 358360 485432
rect 239732 485392 239738 485404
rect 358354 485392 358360 485404
rect 358412 485392 358418 485444
rect 64138 485324 64144 485376
rect 64196 485364 64202 485376
rect 72418 485364 72424 485376
rect 64196 485336 72424 485364
rect 64196 485324 64202 485336
rect 72418 485324 72424 485336
rect 72476 485324 72482 485376
rect 73890 485324 73896 485376
rect 73948 485364 73954 485376
rect 106366 485364 106372 485376
rect 73948 485336 106372 485364
rect 73948 485324 73954 485336
rect 106366 485324 106372 485336
rect 106424 485324 106430 485376
rect 186314 485324 186320 485376
rect 186372 485364 186378 485376
rect 193858 485364 193864 485376
rect 186372 485336 193864 485364
rect 186372 485324 186378 485336
rect 193858 485324 193864 485336
rect 193916 485324 193922 485376
rect 208946 485324 208952 485376
rect 209004 485364 209010 485376
rect 218146 485364 218152 485376
rect 209004 485336 218152 485364
rect 209004 485324 209010 485336
rect 218146 485324 218152 485336
rect 218204 485324 218210 485376
rect 234522 485324 234528 485376
rect 234580 485364 234586 485376
rect 363598 485364 363604 485376
rect 234580 485336 363604 485364
rect 234580 485324 234586 485336
rect 363598 485324 363604 485336
rect 363656 485324 363662 485376
rect 54662 485256 54668 485308
rect 54720 485296 54726 485308
rect 102410 485296 102416 485308
rect 54720 485268 102416 485296
rect 54720 485256 54726 485268
rect 102410 485256 102416 485268
rect 102468 485256 102474 485308
rect 148226 485256 148232 485308
rect 148284 485296 148290 485308
rect 148284 485268 186452 485296
rect 148284 485256 148290 485268
rect 51810 485188 51816 485240
rect 51868 485228 51874 485240
rect 99742 485228 99748 485240
rect 51868 485200 99748 485228
rect 51868 485188 51874 485200
rect 99742 485188 99748 485200
rect 99800 485188 99806 485240
rect 139210 485188 139216 485240
rect 139268 485228 139274 485240
rect 186314 485228 186320 485240
rect 139268 485200 186320 485228
rect 139268 485188 139274 485200
rect 186314 485188 186320 485200
rect 186372 485188 186378 485240
rect 186424 485228 186452 485268
rect 195238 485256 195244 485308
rect 195296 485296 195302 485308
rect 199378 485296 199384 485308
rect 195296 485268 199384 485296
rect 195296 485256 195302 485268
rect 199378 485256 199384 485268
rect 199436 485256 199442 485308
rect 217410 485296 217416 485308
rect 205606 485268 217416 485296
rect 197354 485228 197360 485240
rect 186424 485200 197360 485228
rect 197354 485188 197360 485200
rect 197412 485188 197418 485240
rect 199838 485188 199844 485240
rect 199896 485228 199902 485240
rect 205606 485228 205634 485268
rect 217410 485256 217416 485268
rect 217468 485256 217474 485308
rect 233234 485256 233240 485308
rect 233292 485296 233298 485308
rect 366450 485296 366456 485308
rect 233292 485268 366456 485296
rect 233292 485256 233298 485268
rect 366450 485256 366456 485268
rect 366508 485256 366514 485308
rect 219158 485228 219164 485240
rect 199896 485200 205634 485228
rect 215266 485200 219164 485228
rect 199896 485188 199902 485200
rect 45462 485120 45468 485172
rect 45520 485160 45526 485172
rect 105538 485160 105544 485172
rect 45520 485132 105544 485160
rect 45520 485120 45526 485132
rect 105538 485120 105544 485132
rect 105596 485120 105602 485172
rect 110322 485120 110328 485172
rect 110380 485160 110386 485172
rect 164878 485160 164884 485172
rect 110380 485132 164884 485160
rect 110380 485120 110386 485132
rect 164878 485120 164884 485132
rect 164936 485120 164942 485172
rect 166258 485120 166264 485172
rect 166316 485160 166322 485172
rect 202230 485160 202236 485172
rect 166316 485132 202236 485160
rect 166316 485120 166322 485132
rect 202230 485120 202236 485132
rect 202288 485120 202294 485172
rect 205450 485120 205456 485172
rect 205508 485160 205514 485172
rect 215266 485160 215294 485200
rect 219158 485188 219164 485200
rect 219216 485188 219222 485240
rect 225598 485188 225604 485240
rect 225656 485228 225662 485240
rect 358170 485228 358176 485240
rect 225656 485200 358176 485228
rect 225656 485188 225662 485200
rect 358170 485188 358176 485200
rect 358228 485188 358234 485240
rect 205508 485132 215294 485160
rect 205508 485120 205514 485132
rect 219066 485120 219072 485172
rect 219124 485160 219130 485172
rect 219710 485160 219716 485172
rect 219124 485132 219716 485160
rect 219124 485120 219130 485132
rect 219710 485120 219716 485132
rect 219768 485120 219774 485172
rect 224034 485120 224040 485172
rect 224092 485160 224098 485172
rect 360838 485160 360844 485172
rect 224092 485132 360844 485160
rect 224092 485120 224098 485132
rect 360838 485120 360844 485132
rect 360896 485120 360902 485172
rect 56226 485052 56232 485104
rect 56284 485092 56290 485104
rect 90542 485092 90548 485104
rect 56284 485064 90548 485092
rect 56284 485052 56290 485064
rect 90542 485052 90548 485064
rect 90600 485052 90606 485104
rect 95418 485052 95424 485104
rect 95476 485092 95482 485104
rect 167822 485092 167828 485104
rect 95476 485064 167828 485092
rect 95476 485052 95482 485064
rect 167822 485052 167828 485064
rect 167880 485052 167886 485104
rect 182266 485052 182272 485104
rect 182324 485092 182330 485104
rect 208394 485092 208400 485104
rect 182324 485064 208400 485092
rect 182324 485052 182330 485064
rect 208394 485052 208400 485064
rect 208452 485052 208458 485104
rect 209498 485052 209504 485104
rect 209556 485092 209562 485104
rect 221734 485092 221740 485104
rect 209556 485064 221740 485092
rect 209556 485052 209562 485064
rect 221734 485052 221740 485064
rect 221792 485052 221798 485104
rect 223482 485052 223488 485104
rect 223540 485092 223546 485104
rect 371878 485092 371884 485104
rect 223540 485064 371884 485092
rect 223540 485052 223546 485064
rect 371878 485052 371884 485064
rect 371936 485052 371942 485104
rect 58618 484984 58624 485036
rect 58676 485024 58682 485036
rect 81250 485024 81256 485036
rect 58676 484996 81256 485024
rect 58676 484984 58682 484996
rect 81250 484984 81256 484996
rect 81308 484984 81314 485036
rect 149882 484984 149888 485036
rect 149940 485024 149946 485036
rect 197354 485024 197360 485036
rect 149940 484996 197360 485024
rect 149940 484984 149946 484996
rect 197354 484984 197360 484996
rect 197412 484984 197418 485036
rect 202690 484984 202696 485036
rect 202748 485024 202754 485036
rect 210142 485024 210148 485036
rect 202748 484996 210148 485024
rect 202748 484984 202754 484996
rect 210142 484984 210148 484996
rect 210200 484984 210206 485036
rect 53650 484916 53656 484968
rect 53708 484956 53714 484968
rect 74442 484956 74448 484968
rect 53708 484928 74448 484956
rect 53708 484916 53714 484928
rect 74442 484916 74448 484928
rect 74500 484916 74506 484968
rect 156598 484916 156604 484968
rect 156656 484956 156662 484968
rect 166166 484956 166172 484968
rect 156656 484928 166172 484956
rect 156656 484916 156662 484928
rect 166166 484916 166172 484928
rect 166224 484916 166230 484968
rect 166258 484916 166264 484968
rect 166316 484956 166322 484968
rect 201494 484956 201500 484968
rect 166316 484928 201500 484956
rect 166316 484916 166322 484928
rect 201494 484916 201500 484928
rect 201552 484916 201558 484968
rect 209038 484916 209044 484968
rect 209096 484956 209102 484968
rect 219158 484956 219164 484968
rect 209096 484928 219164 484956
rect 209096 484916 209102 484928
rect 219158 484916 219164 484928
rect 219216 484916 219222 484968
rect 59170 484848 59176 484900
rect 59228 484888 59234 484900
rect 69658 484888 69664 484900
rect 59228 484860 69664 484888
rect 59228 484848 59234 484860
rect 69658 484848 69664 484860
rect 69716 484848 69722 484900
rect 84378 484888 84384 484900
rect 69876 484860 84384 484888
rect 53282 484780 53288 484832
rect 53340 484820 53346 484832
rect 53340 484792 64874 484820
rect 53340 484780 53346 484792
rect 64846 484684 64874 484792
rect 68278 484712 68284 484764
rect 68336 484752 68342 484764
rect 69876 484752 69904 484860
rect 84378 484848 84384 484860
rect 84436 484848 84442 484900
rect 139394 484848 139400 484900
rect 139452 484888 139458 484900
rect 185578 484888 185584 484900
rect 139452 484860 185584 484888
rect 139452 484848 139458 484860
rect 185578 484848 185584 484860
rect 185636 484848 185642 484900
rect 191190 484848 191196 484900
rect 191248 484888 191254 484900
rect 200482 484888 200488 484900
rect 191248 484860 200488 484888
rect 191248 484848 191254 484860
rect 200482 484848 200488 484860
rect 200540 484848 200546 484900
rect 157426 484780 157432 484832
rect 157484 484820 157490 484832
rect 208394 484820 208400 484832
rect 157484 484792 208400 484820
rect 157484 484780 157490 484792
rect 208394 484780 208400 484792
rect 208452 484780 208458 484832
rect 68336 484724 69904 484752
rect 68336 484712 68342 484724
rect 155586 484712 155592 484764
rect 155644 484752 155650 484764
rect 166258 484752 166264 484764
rect 155644 484724 166264 484752
rect 155644 484712 155650 484724
rect 166258 484712 166264 484724
rect 166316 484712 166322 484764
rect 167822 484712 167828 484764
rect 167880 484752 167886 484764
rect 182818 484752 182824 484764
rect 167880 484724 182824 484752
rect 167880 484712 167886 484724
rect 182818 484712 182824 484724
rect 182876 484712 182882 484764
rect 77754 484684 77760 484696
rect 64846 484656 77760 484684
rect 77754 484644 77760 484656
rect 77812 484644 77818 484696
rect 195146 484372 195152 484424
rect 195204 484412 195210 484424
rect 197078 484412 197084 484424
rect 195204 484384 197084 484412
rect 195204 484372 195210 484384
rect 197078 484372 197084 484384
rect 197136 484372 197142 484424
rect 213362 484372 213368 484424
rect 213420 484412 213426 484424
rect 214926 484412 214932 484424
rect 213420 484384 214932 484412
rect 213420 484372 213426 484384
rect 214926 484372 214932 484384
rect 214984 484372 214990 484424
rect 219986 484372 219992 484424
rect 220044 484412 220050 484424
rect 222654 484412 222660 484424
rect 220044 484384 222660 484412
rect 220044 484372 220050 484384
rect 222654 484372 222660 484384
rect 222712 484372 222718 484424
rect 203702 484304 203708 484356
rect 203760 484344 203766 484356
rect 209590 484344 209596 484356
rect 203760 484316 209596 484344
rect 203760 484304 203766 484316
rect 209590 484304 209596 484316
rect 209648 484304 209654 484356
rect 161566 484236 161572 484288
rect 161624 484276 161630 484288
rect 162762 484276 162768 484288
rect 161624 484248 162768 484276
rect 161624 484236 161630 484248
rect 162762 484236 162768 484248
rect 162820 484236 162826 484288
rect 226610 484236 226616 484288
rect 226668 484276 226674 484288
rect 227622 484276 227628 484288
rect 226668 484248 227628 484276
rect 226668 484236 226674 484248
rect 227622 484236 227628 484248
rect 227680 484236 227686 484288
rect 92566 484168 92572 484220
rect 92624 484208 92630 484220
rect 93302 484208 93308 484220
rect 92624 484180 93308 484208
rect 92624 484168 92630 484180
rect 93302 484168 93308 484180
rect 93360 484168 93366 484220
rect 103514 484168 103520 484220
rect 103572 484208 103578 484220
rect 104342 484208 104348 484220
rect 103572 484180 104348 484208
rect 103572 484168 103578 484180
rect 104342 484168 104348 484180
rect 104400 484168 104406 484220
rect 129826 484168 129832 484220
rect 129884 484208 129890 484220
rect 130654 484208 130660 484220
rect 129884 484180 130660 484208
rect 129884 484168 129890 484180
rect 130654 484168 130660 484180
rect 130712 484168 130718 484220
rect 143626 484168 143632 484220
rect 143684 484208 143690 484220
rect 143902 484208 143908 484220
rect 143684 484180 143908 484208
rect 143684 484168 143690 484180
rect 143902 484168 143908 484180
rect 143960 484168 143966 484220
rect 161474 484168 161480 484220
rect 161532 484208 161538 484220
rect 161934 484208 161940 484220
rect 161532 484180 161940 484208
rect 161532 484168 161538 484180
rect 161934 484168 161940 484180
rect 161992 484168 161998 484220
rect 219526 484168 219532 484220
rect 219584 484208 219590 484220
rect 219894 484208 219900 484220
rect 219584 484180 219900 484208
rect 219584 484168 219590 484180
rect 219894 484168 219900 484180
rect 219952 484168 219958 484220
rect 265158 484168 265164 484220
rect 265216 484208 265222 484220
rect 265894 484208 265900 484220
rect 265216 484180 265900 484208
rect 265216 484168 265222 484180
rect 265894 484168 265900 484180
rect 265952 484168 265958 484220
rect 266446 484168 266452 484220
rect 266504 484208 266510 484220
rect 267182 484208 267188 484220
rect 266504 484180 267188 484208
rect 266504 484168 266510 484180
rect 267182 484168 267188 484180
rect 267240 484168 267246 484220
rect 60734 484100 60740 484152
rect 60792 484140 60798 484152
rect 61102 484140 61108 484152
rect 60792 484112 61108 484140
rect 60792 484100 60798 484112
rect 61102 484100 61108 484112
rect 61160 484100 61166 484152
rect 62114 484100 62120 484152
rect 62172 484140 62178 484152
rect 62942 484140 62948 484152
rect 62172 484112 62948 484140
rect 62172 484100 62178 484112
rect 62942 484100 62948 484112
rect 63000 484100 63006 484152
rect 64874 484100 64880 484152
rect 64932 484140 64938 484152
rect 65518 484140 65524 484152
rect 64932 484112 65524 484140
rect 64932 484100 64938 484112
rect 65518 484100 65524 484112
rect 65576 484100 65582 484152
rect 67726 484100 67732 484152
rect 67784 484140 67790 484152
rect 68186 484140 68192 484152
rect 67784 484112 68192 484140
rect 67784 484100 67790 484112
rect 68186 484100 68192 484112
rect 68244 484100 68250 484152
rect 69014 484100 69020 484152
rect 69072 484140 69078 484152
rect 69566 484140 69572 484152
rect 69072 484112 69572 484140
rect 69072 484100 69078 484112
rect 69566 484100 69572 484112
rect 69624 484100 69630 484152
rect 92474 484100 92480 484152
rect 92532 484140 92538 484152
rect 92934 484140 92940 484152
rect 92532 484112 92940 484140
rect 92532 484100 92538 484112
rect 92934 484100 92940 484112
rect 92992 484100 92998 484152
rect 93854 484100 93860 484152
rect 93912 484140 93918 484152
rect 94590 484140 94596 484152
rect 93912 484112 94596 484140
rect 93912 484100 93918 484112
rect 94590 484100 94596 484112
rect 94648 484100 94654 484152
rect 99466 484100 99472 484152
rect 99524 484140 99530 484152
rect 100294 484140 100300 484152
rect 99524 484112 100300 484140
rect 99524 484100 99530 484112
rect 100294 484100 100300 484112
rect 100352 484100 100358 484152
rect 103606 484100 103612 484152
rect 103664 484140 103670 484152
rect 103790 484140 103796 484152
rect 103664 484112 103796 484140
rect 103664 484100 103670 484112
rect 103790 484100 103796 484112
rect 103848 484100 103854 484152
rect 107654 484100 107660 484152
rect 107712 484140 107718 484152
rect 107838 484140 107844 484152
rect 107712 484112 107844 484140
rect 107712 484100 107718 484112
rect 107838 484100 107844 484112
rect 107896 484100 107902 484152
rect 122834 484100 122840 484152
rect 122892 484140 122898 484152
rect 123662 484140 123668 484152
rect 122892 484112 123668 484140
rect 122892 484100 122898 484112
rect 123662 484100 123668 484112
rect 123720 484100 123726 484152
rect 124306 484100 124312 484152
rect 124364 484140 124370 484152
rect 124950 484140 124956 484152
rect 124364 484112 124956 484140
rect 124364 484100 124370 484112
rect 124950 484100 124956 484112
rect 125008 484100 125014 484152
rect 125594 484100 125600 484152
rect 125652 484140 125658 484152
rect 126330 484140 126336 484152
rect 125652 484112 126336 484140
rect 125652 484100 125658 484112
rect 126330 484100 126336 484112
rect 126388 484100 126394 484152
rect 129918 484100 129924 484152
rect 129976 484140 129982 484152
rect 130286 484140 130292 484152
rect 129976 484112 130292 484140
rect 129976 484100 129982 484112
rect 130286 484100 130292 484112
rect 130344 484100 130350 484152
rect 131114 484100 131120 484152
rect 131172 484140 131178 484152
rect 132126 484140 132132 484152
rect 131172 484112 132132 484140
rect 131172 484100 131178 484112
rect 132126 484100 132132 484112
rect 132184 484100 132190 484152
rect 133874 484100 133880 484152
rect 133932 484140 133938 484152
rect 134334 484140 134340 484152
rect 133932 484112 134340 484140
rect 133932 484100 133938 484112
rect 134334 484100 134340 484112
rect 134392 484100 134398 484152
rect 139394 484100 139400 484152
rect 139452 484140 139458 484152
rect 140038 484140 140044 484152
rect 139452 484112 140044 484140
rect 139452 484100 139458 484112
rect 140038 484100 140044 484112
rect 140096 484100 140102 484152
rect 140866 484100 140872 484152
rect 140924 484140 140930 484152
rect 141694 484140 141700 484152
rect 140924 484112 141700 484140
rect 140924 484100 140930 484112
rect 141694 484100 141700 484112
rect 141752 484100 141758 484152
rect 142154 484100 142160 484152
rect 142212 484140 142218 484152
rect 142614 484140 142620 484152
rect 142212 484112 142620 484140
rect 142212 484100 142218 484112
rect 142614 484100 142620 484112
rect 142672 484100 142678 484152
rect 143534 484100 143540 484152
rect 143592 484140 143598 484152
rect 144454 484140 144460 484152
rect 143592 484112 144460 484140
rect 143592 484100 143598 484112
rect 144454 484100 144460 484112
rect 144512 484100 144518 484152
rect 147674 484100 147680 484152
rect 147732 484140 147738 484152
rect 148318 484140 148324 484152
rect 147732 484112 148324 484140
rect 147732 484100 147738 484112
rect 148318 484100 148324 484112
rect 148376 484100 148382 484152
rect 160094 484100 160100 484152
rect 160152 484140 160158 484152
rect 160646 484140 160652 484152
rect 160152 484112 160652 484140
rect 160152 484100 160158 484112
rect 160646 484100 160652 484112
rect 160704 484100 160710 484152
rect 161566 484100 161572 484152
rect 161624 484140 161630 484152
rect 162486 484140 162492 484152
rect 161624 484112 162492 484140
rect 161624 484100 161630 484112
rect 162486 484100 162492 484112
rect 162544 484100 162550 484152
rect 162854 484100 162860 484152
rect 162912 484140 162918 484152
rect 163774 484140 163780 484152
rect 162912 484112 163780 484140
rect 162912 484100 162918 484112
rect 163774 484100 163780 484112
rect 163832 484100 163838 484152
rect 196710 484100 196716 484152
rect 196768 484140 196774 484152
rect 196894 484140 196900 484152
rect 196768 484112 196900 484140
rect 196768 484100 196774 484112
rect 196894 484100 196900 484112
rect 196952 484100 196958 484152
rect 197446 484100 197452 484152
rect 197504 484140 197510 484152
rect 198366 484140 198372 484152
rect 197504 484112 198372 484140
rect 197504 484100 197510 484112
rect 198366 484100 198372 484112
rect 198424 484100 198430 484152
rect 198734 484100 198740 484152
rect 198792 484140 198798 484152
rect 198918 484140 198924 484152
rect 198792 484112 198924 484140
rect 198792 484100 198798 484112
rect 198918 484100 198924 484112
rect 198976 484100 198982 484152
rect 204438 484100 204444 484152
rect 204496 484140 204502 484152
rect 205174 484140 205180 484152
rect 204496 484112 205180 484140
rect 204496 484100 204502 484112
rect 205174 484100 205180 484112
rect 205232 484100 205238 484152
rect 215386 484100 215392 484152
rect 215444 484140 215450 484152
rect 216214 484140 216220 484152
rect 215444 484112 216220 484140
rect 215444 484100 215450 484112
rect 216214 484100 216220 484112
rect 216272 484100 216278 484152
rect 216766 484100 216772 484152
rect 216824 484140 216830 484152
rect 217502 484140 217508 484152
rect 216824 484112 217508 484140
rect 216824 484100 216830 484112
rect 217502 484100 217508 484112
rect 217560 484100 217566 484152
rect 219618 484100 219624 484152
rect 219676 484140 219682 484152
rect 220078 484140 220084 484152
rect 219676 484112 220084 484140
rect 219676 484100 219682 484112
rect 220078 484100 220084 484112
rect 220136 484100 220142 484152
rect 227714 484100 227720 484152
rect 227772 484140 227778 484152
rect 228542 484140 228548 484152
rect 227772 484112 228548 484140
rect 227772 484100 227778 484112
rect 228542 484100 228548 484112
rect 228600 484100 228606 484152
rect 229094 484100 229100 484152
rect 229152 484140 229158 484152
rect 229462 484140 229468 484152
rect 229152 484112 229468 484140
rect 229152 484100 229158 484112
rect 229462 484100 229468 484112
rect 229520 484100 229526 484152
rect 235994 484100 236000 484152
rect 236052 484140 236058 484152
rect 236822 484140 236828 484152
rect 236052 484112 236828 484140
rect 236052 484100 236058 484112
rect 236822 484100 236828 484112
rect 236880 484100 236886 484152
rect 241514 484100 241520 484152
rect 241572 484140 241578 484152
rect 242158 484140 242164 484152
rect 241572 484112 242164 484140
rect 241572 484100 241578 484112
rect 242158 484100 242164 484112
rect 242216 484100 242222 484152
rect 265066 484100 265072 484152
rect 265124 484140 265130 484152
rect 265526 484140 265532 484152
rect 265124 484112 265532 484140
rect 265124 484100 265130 484112
rect 265526 484100 265532 484112
rect 265584 484100 265590 484152
rect 266354 484100 266360 484152
rect 266412 484140 266418 484152
rect 266814 484140 266820 484152
rect 266412 484112 266820 484140
rect 266412 484100 266418 484112
rect 266814 484100 266820 484112
rect 266872 484100 266878 484152
rect 284294 484100 284300 484152
rect 284352 484140 284358 484152
rect 284846 484140 284852 484152
rect 284352 484112 284852 484140
rect 284352 484100 284358 484112
rect 284846 484100 284852 484112
rect 284904 484100 284910 484152
rect 287054 484100 287060 484152
rect 287112 484140 287118 484152
rect 287974 484140 287980 484152
rect 287112 484112 287980 484140
rect 287112 484100 287118 484112
rect 287974 484100 287980 484112
rect 288032 484100 288038 484152
rect 289906 484100 289912 484152
rect 289964 484140 289970 484152
rect 290550 484140 290556 484152
rect 289964 484112 290556 484140
rect 289964 484100 289970 484112
rect 290550 484100 290556 484112
rect 290608 484100 290614 484152
rect 291286 484100 291292 484152
rect 291344 484140 291350 484152
rect 291930 484140 291936 484152
rect 291344 484112 291936 484140
rect 291344 484100 291350 484112
rect 291930 484100 291936 484112
rect 291988 484100 291994 484152
rect 264974 484032 264980 484084
rect 265032 484072 265038 484084
rect 265342 484072 265348 484084
rect 265032 484044 265348 484072
rect 265032 484032 265038 484044
rect 265342 484032 265348 484044
rect 265400 484032 265406 484084
rect 281442 484032 281448 484084
rect 281500 484072 281506 484084
rect 281500 484044 284708 484072
rect 281500 484032 281506 484044
rect 60826 483964 60832 484016
rect 60884 484004 60890 484016
rect 61654 484004 61660 484016
rect 60884 483976 61660 484004
rect 60884 483964 60890 483976
rect 61654 483964 61660 483976
rect 61712 483964 61718 484016
rect 284680 484004 284708 484044
rect 286962 484032 286968 484084
rect 287020 484072 287026 484084
rect 356882 484072 356888 484084
rect 287020 484044 356888 484072
rect 287020 484032 287026 484044
rect 356882 484032 356888 484044
rect 356940 484032 356946 484084
rect 376386 484004 376392 484016
rect 284680 483976 376392 484004
rect 376386 483964 376392 483976
rect 376444 483964 376450 484016
rect 269022 483896 269028 483948
rect 269080 483936 269086 483948
rect 370406 483936 370412 483948
rect 269080 483908 370412 483936
rect 269080 483896 269086 483908
rect 370406 483896 370412 483908
rect 370464 483896 370470 483948
rect 268010 483828 268016 483880
rect 268068 483868 268074 483880
rect 377306 483868 377312 483880
rect 268068 483840 377312 483868
rect 268068 483828 268074 483840
rect 377306 483828 377312 483840
rect 377364 483828 377370 483880
rect 177298 483760 177304 483812
rect 177356 483800 177362 483812
rect 205174 483800 205180 483812
rect 177356 483772 205180 483800
rect 177356 483760 177362 483772
rect 205174 483760 205180 483772
rect 205232 483760 205238 483812
rect 246022 483760 246028 483812
rect 246080 483800 246086 483812
rect 369210 483800 369216 483812
rect 246080 483772 369216 483800
rect 246080 483760 246086 483772
rect 369210 483760 369216 483772
rect 369268 483760 369274 483812
rect 60642 483692 60648 483744
rect 60700 483732 60706 483744
rect 80698 483732 80704 483744
rect 60700 483704 80704 483732
rect 60700 483692 60706 483704
rect 80698 483692 80704 483704
rect 80756 483692 80762 483744
rect 162762 483692 162768 483744
rect 162820 483732 162826 483744
rect 215938 483732 215944 483744
rect 162820 483704 215944 483732
rect 162820 483692 162826 483704
rect 215938 483692 215944 483704
rect 215996 483692 216002 483744
rect 227898 483692 227904 483744
rect 227956 483732 227962 483744
rect 362218 483732 362224 483744
rect 227956 483704 362224 483732
rect 227956 483692 227962 483704
rect 362218 483692 362224 483704
rect 362276 483692 362282 483744
rect 56778 483624 56784 483676
rect 56836 483664 56842 483676
rect 113450 483664 113456 483676
rect 56836 483636 113456 483664
rect 56836 483624 56842 483636
rect 113450 483624 113456 483636
rect 113508 483624 113514 483676
rect 160002 483624 160008 483676
rect 160060 483664 160066 483676
rect 214558 483664 214564 483676
rect 160060 483636 214564 483664
rect 160060 483624 160066 483636
rect 214558 483624 214564 483636
rect 214616 483624 214622 483676
rect 227622 483624 227628 483676
rect 227680 483664 227686 483676
rect 370498 483664 370504 483676
rect 227680 483636 370504 483664
rect 227680 483624 227686 483636
rect 370498 483624 370504 483636
rect 370556 483624 370562 483676
rect 201494 483488 201500 483540
rect 201552 483528 201558 483540
rect 201678 483528 201684 483540
rect 201552 483500 201684 483528
rect 201552 483488 201558 483500
rect 201678 483488 201684 483500
rect 201736 483488 201742 483540
rect 223574 483352 223580 483404
rect 223632 483392 223638 483404
rect 224126 483392 224132 483404
rect 223632 483364 224132 483392
rect 223632 483352 223638 483364
rect 224126 483352 224132 483364
rect 224184 483352 224190 483404
rect 50430 482944 50436 482996
rect 50488 482984 50494 482996
rect 97166 482984 97172 482996
rect 50488 482956 97172 482984
rect 50488 482944 50494 482956
rect 97166 482944 97172 482956
rect 97224 482944 97230 482996
rect 50522 482876 50528 482928
rect 50580 482916 50586 482928
rect 98454 482916 98460 482928
rect 50580 482888 98460 482916
rect 50580 482876 50586 482888
rect 98454 482876 98460 482888
rect 98512 482876 98518 482928
rect 299382 482876 299388 482928
rect 299440 482916 299446 482928
rect 364058 482916 364064 482928
rect 299440 482888 364064 482916
rect 299440 482876 299446 482888
rect 364058 482876 364064 482888
rect 364116 482876 364122 482928
rect 48038 482808 48044 482860
rect 48096 482848 48102 482860
rect 97994 482848 98000 482860
rect 48096 482820 98000 482848
rect 48096 482808 48102 482820
rect 97994 482808 98000 482820
rect 98052 482808 98058 482860
rect 284754 482808 284760 482860
rect 284812 482848 284818 482860
rect 359826 482848 359832 482860
rect 284812 482820 359832 482848
rect 284812 482808 284818 482820
rect 359826 482808 359832 482820
rect 359884 482808 359890 482860
rect 48130 482740 48136 482792
rect 48188 482780 48194 482792
rect 111702 482780 111708 482792
rect 48188 482752 111708 482780
rect 48188 482740 48194 482752
rect 111702 482740 111708 482752
rect 111760 482740 111766 482792
rect 177114 482740 177120 482792
rect 177172 482780 177178 482792
rect 203610 482780 203616 482792
rect 177172 482752 203616 482780
rect 177172 482740 177178 482752
rect 203610 482740 203616 482752
rect 203668 482740 203674 482792
rect 280062 482740 280068 482792
rect 280120 482780 280126 482792
rect 361298 482780 361304 482792
rect 280120 482752 361304 482780
rect 280120 482740 280126 482752
rect 361298 482740 361304 482752
rect 361356 482740 361362 482792
rect 46658 482672 46664 482724
rect 46716 482712 46722 482724
rect 111242 482712 111248 482724
rect 46716 482684 111248 482712
rect 46716 482672 46722 482684
rect 111242 482672 111248 482684
rect 111300 482672 111306 482724
rect 173434 482672 173440 482724
rect 173492 482712 173498 482724
rect 216030 482712 216036 482724
rect 173492 482684 216036 482712
rect 173492 482672 173498 482684
rect 216030 482672 216036 482684
rect 216088 482672 216094 482724
rect 278682 482672 278688 482724
rect 278740 482712 278746 482724
rect 362678 482712 362684 482724
rect 278740 482684 362684 482712
rect 278740 482672 278746 482684
rect 362678 482672 362684 482684
rect 362736 482672 362742 482724
rect 50614 482604 50620 482656
rect 50672 482644 50678 482656
rect 115658 482644 115664 482656
rect 50672 482616 115664 482644
rect 50672 482604 50678 482616
rect 115658 482604 115664 482616
rect 115716 482604 115722 482656
rect 138474 482604 138480 482656
rect 138532 482644 138538 482656
rect 138532 482616 142154 482644
rect 138532 482604 138538 482616
rect 46382 482536 46388 482588
rect 46440 482576 46446 482588
rect 112070 482576 112076 482588
rect 46440 482548 112076 482576
rect 46440 482536 46446 482548
rect 112070 482536 112076 482548
rect 112128 482536 112134 482588
rect 140774 482536 140780 482588
rect 140832 482576 140838 482588
rect 141326 482576 141332 482588
rect 140832 482548 141332 482576
rect 140832 482536 140838 482548
rect 141326 482536 141332 482548
rect 141384 482536 141390 482588
rect 142126 482576 142154 482616
rect 165522 482604 165528 482656
rect 165580 482644 165586 482656
rect 214650 482644 214656 482656
rect 165580 482616 214656 482644
rect 165580 482604 165586 482616
rect 214650 482604 214656 482616
rect 214708 482604 214714 482656
rect 272426 482604 272432 482656
rect 272484 482644 272490 482656
rect 369670 482644 369676 482656
rect 272484 482616 369676 482644
rect 272484 482604 272490 482616
rect 369670 482604 369676 482616
rect 369728 482604 369734 482656
rect 197170 482576 197176 482588
rect 142126 482548 197176 482576
rect 197170 482536 197176 482548
rect 197228 482536 197234 482588
rect 242894 482536 242900 482588
rect 242952 482576 242958 482588
rect 243078 482576 243084 482588
rect 242952 482548 243084 482576
rect 242952 482536 242958 482548
rect 243078 482536 243084 482548
rect 243136 482536 243142 482588
rect 257522 482536 257528 482588
rect 257580 482576 257586 482588
rect 362494 482576 362500 482588
rect 257580 482548 362500 482576
rect 257580 482536 257586 482548
rect 362494 482536 362500 482548
rect 362552 482536 362558 482588
rect 49050 482468 49056 482520
rect 49108 482508 49114 482520
rect 115198 482508 115204 482520
rect 49108 482480 115204 482508
rect 49108 482468 49114 482480
rect 115198 482468 115204 482480
rect 115256 482468 115262 482520
rect 135714 482468 135720 482520
rect 135772 482508 135778 482520
rect 197906 482508 197912 482520
rect 135772 482480 197912 482508
rect 135772 482468 135778 482480
rect 197906 482468 197912 482480
rect 197964 482468 197970 482520
rect 261386 482468 261392 482520
rect 261444 482508 261450 482520
rect 369486 482508 369492 482520
rect 261444 482480 369492 482508
rect 261444 482468 261450 482480
rect 369486 482468 369492 482480
rect 369544 482468 369550 482520
rect 46290 482400 46296 482452
rect 46348 482440 46354 482452
rect 112530 482440 112536 482452
rect 46348 482412 112536 482440
rect 46348 482400 46354 482412
rect 112530 482400 112536 482412
rect 112588 482400 112594 482452
rect 138842 482400 138848 482452
rect 138900 482440 138906 482452
rect 201770 482440 201776 482452
rect 138900 482412 201776 482440
rect 138900 482400 138906 482412
rect 201770 482400 201776 482412
rect 201828 482400 201834 482452
rect 255222 482400 255228 482452
rect 255280 482440 255286 482452
rect 369578 482440 369584 482452
rect 255280 482412 369584 482440
rect 255280 482400 255286 482412
rect 369578 482400 369584 482412
rect 369636 482400 369642 482452
rect 46750 482332 46756 482384
rect 46808 482372 46814 482384
rect 119614 482372 119620 482384
rect 46808 482344 119620 482372
rect 46808 482332 46814 482344
rect 119614 482332 119620 482344
rect 119672 482332 119678 482384
rect 137922 482332 137928 482384
rect 137980 482372 137986 482384
rect 203150 482372 203156 482384
rect 137980 482344 203156 482372
rect 137980 482332 137986 482344
rect 203150 482332 203156 482344
rect 203208 482332 203214 482384
rect 244642 482332 244648 482384
rect 244700 482372 244706 482384
rect 372062 482372 372068 482384
rect 244700 482344 372068 482372
rect 244700 482332 244706 482344
rect 372062 482332 372068 482344
rect 372120 482332 372126 482384
rect 57238 482264 57244 482316
rect 57296 482304 57302 482316
rect 135898 482304 135904 482316
rect 57296 482276 135904 482304
rect 57296 482264 57302 482276
rect 135898 482264 135904 482276
rect 135956 482264 135962 482316
rect 137554 482264 137560 482316
rect 137612 482304 137618 482316
rect 204622 482304 204628 482316
rect 137612 482276 204628 482304
rect 137612 482264 137618 482276
rect 204622 482264 204628 482276
rect 204680 482264 204686 482316
rect 248322 482264 248328 482316
rect 248380 482304 248386 482316
rect 378778 482304 378784 482316
rect 248380 482276 378784 482304
rect 248380 482264 248386 482276
rect 378778 482264 378784 482276
rect 378836 482264 378842 482316
rect 51626 482196 51632 482248
rect 51684 482236 51690 482248
rect 97534 482236 97540 482248
rect 51684 482208 97540 482236
rect 51684 482196 51690 482208
rect 97534 482196 97540 482208
rect 97592 482196 97598 482248
rect 54570 482128 54576 482180
rect 54628 482168 54634 482180
rect 96706 482168 96712 482180
rect 54628 482140 96712 482168
rect 54628 482128 54634 482140
rect 96706 482128 96712 482140
rect 96764 482128 96770 482180
rect 58802 482060 58808 482112
rect 58860 482100 58866 482112
rect 96246 482100 96252 482112
rect 58860 482072 96252 482100
rect 58860 482060 58866 482072
rect 96246 482060 96252 482072
rect 96304 482060 96310 482112
rect 125686 481992 125692 482044
rect 125744 482032 125750 482044
rect 125870 482032 125876 482044
rect 125744 482004 125876 482032
rect 125744 481992 125750 482004
rect 125870 481992 125876 482004
rect 125928 481992 125934 482044
rect 289722 481312 289728 481364
rect 289780 481352 289786 481364
rect 372430 481352 372436 481364
rect 289780 481324 372436 481352
rect 289780 481312 289786 481324
rect 372430 481312 372436 481324
rect 372488 481312 372494 481364
rect 270034 481244 270040 481296
rect 270092 481284 270098 481296
rect 358630 481284 358636 481296
rect 270092 481256 358636 481284
rect 270092 481244 270098 481256
rect 358630 481244 358636 481256
rect 358688 481244 358694 481296
rect 262214 481176 262220 481228
rect 262272 481216 262278 481228
rect 262582 481216 262588 481228
rect 262272 481188 262588 481216
rect 262272 481176 262278 481188
rect 262582 481176 262588 481188
rect 262640 481176 262646 481228
rect 270402 481176 270408 481228
rect 270460 481216 270466 481228
rect 359458 481216 359464 481228
rect 270460 481188 359464 481216
rect 270460 481176 270466 481188
rect 359458 481176 359464 481188
rect 359516 481176 359522 481228
rect 189166 481108 189172 481160
rect 189224 481148 189230 481160
rect 189350 481148 189356 481160
rect 189224 481120 189356 481148
rect 189224 481108 189230 481120
rect 189350 481108 189356 481120
rect 189408 481108 189414 481160
rect 251358 481108 251364 481160
rect 251416 481148 251422 481160
rect 251542 481148 251548 481160
rect 251416 481120 251548 481148
rect 251416 481108 251422 481120
rect 251542 481108 251548 481120
rect 251600 481108 251606 481160
rect 271782 481108 271788 481160
rect 271840 481148 271846 481160
rect 377214 481148 377220 481160
rect 271840 481120 377220 481148
rect 271840 481108 271846 481120
rect 377214 481108 377220 481120
rect 377272 481108 377278 481160
rect 74718 481040 74724 481092
rect 74776 481080 74782 481092
rect 74902 481080 74908 481092
rect 74776 481052 74908 481080
rect 74776 481040 74782 481052
rect 74902 481040 74908 481052
rect 74960 481040 74966 481092
rect 168558 481040 168564 481092
rect 168616 481080 168622 481092
rect 168742 481080 168748 481092
rect 168616 481052 168748 481080
rect 168616 481040 168622 481052
rect 168742 481040 168748 481052
rect 168800 481040 168806 481092
rect 176010 481040 176016 481092
rect 176068 481080 176074 481092
rect 209222 481080 209228 481092
rect 176068 481052 209228 481080
rect 176068 481040 176074 481052
rect 209222 481040 209228 481052
rect 209280 481040 209286 481092
rect 212718 481040 212724 481092
rect 212776 481080 212782 481092
rect 212902 481080 212908 481092
rect 212776 481052 212908 481080
rect 212776 481040 212782 481052
rect 212902 481040 212908 481052
rect 212960 481040 212966 481092
rect 244090 481040 244096 481092
rect 244148 481080 244154 481092
rect 363690 481080 363696 481092
rect 244148 481052 363696 481080
rect 244148 481040 244154 481052
rect 363690 481040 363696 481052
rect 363748 481040 363754 481092
rect 57790 480972 57796 481024
rect 57848 481012 57854 481024
rect 114278 481012 114284 481024
rect 57848 480984 114284 481012
rect 57848 480972 57854 480984
rect 114278 480972 114284 480984
rect 114336 480972 114342 481024
rect 160554 480972 160560 481024
rect 160612 481012 160618 481024
rect 211798 481012 211804 481024
rect 160612 480984 211804 481012
rect 160612 480972 160618 480984
rect 211798 480972 211804 480984
rect 211856 480972 211862 481024
rect 253106 480972 253112 481024
rect 253164 481012 253170 481024
rect 374822 481012 374828 481024
rect 253164 480984 374828 481012
rect 253164 480972 253170 480984
rect 374822 480972 374828 480984
rect 374880 480972 374886 481024
rect 3694 480904 3700 480956
rect 3752 480944 3758 480956
rect 434898 480944 434904 480956
rect 3752 480916 434904 480944
rect 3752 480904 3758 480916
rect 434898 480904 434904 480916
rect 434956 480904 434962 480956
rect 70394 480836 70400 480888
rect 70452 480876 70458 480888
rect 70854 480876 70860 480888
rect 70452 480848 70860 480876
rect 70452 480836 70458 480848
rect 70854 480836 70860 480848
rect 70912 480836 70918 480888
rect 74626 480836 74632 480888
rect 74684 480876 74690 480888
rect 75270 480876 75276 480888
rect 74684 480848 75276 480876
rect 74684 480836 74690 480848
rect 75270 480836 75276 480848
rect 75328 480836 75334 480888
rect 75914 480836 75920 480888
rect 75972 480876 75978 480888
rect 76558 480876 76564 480888
rect 75972 480848 76564 480876
rect 75972 480836 75978 480848
rect 76558 480836 76564 480848
rect 76616 480836 76622 480888
rect 81526 480836 81532 480888
rect 81584 480876 81590 480888
rect 82262 480876 82268 480888
rect 81584 480848 82268 480876
rect 81584 480836 81590 480848
rect 82262 480836 82268 480848
rect 82320 480836 82326 480888
rect 82906 480836 82912 480888
rect 82964 480876 82970 480888
rect 83550 480876 83556 480888
rect 82964 480848 83556 480876
rect 82964 480836 82970 480848
rect 83550 480836 83556 480848
rect 83608 480836 83614 480888
rect 84286 480836 84292 480888
rect 84344 480876 84350 480888
rect 84930 480876 84936 480888
rect 84344 480848 84936 480876
rect 84344 480836 84350 480848
rect 84930 480836 84936 480848
rect 84988 480836 84994 480888
rect 86954 480836 86960 480888
rect 87012 480876 87018 480888
rect 87598 480876 87604 480888
rect 87012 480848 87604 480876
rect 87012 480836 87018 480848
rect 87598 480836 87604 480848
rect 87656 480836 87662 480888
rect 88426 480836 88432 480888
rect 88484 480876 88490 480888
rect 89254 480876 89260 480888
rect 88484 480848 89260 480876
rect 88484 480836 88490 480848
rect 89254 480836 89260 480848
rect 89312 480836 89318 480888
rect 167086 480836 167092 480888
rect 167144 480876 167150 480888
rect 167730 480876 167736 480888
rect 167144 480848 167736 480876
rect 167144 480836 167150 480848
rect 167730 480836 167736 480848
rect 167788 480836 167794 480888
rect 168374 480836 168380 480888
rect 168432 480876 168438 480888
rect 169110 480876 169116 480888
rect 168432 480848 169116 480876
rect 168432 480836 168438 480848
rect 169110 480836 169116 480848
rect 169168 480836 169174 480888
rect 169754 480836 169760 480888
rect 169812 480876 169818 480888
rect 170030 480876 170036 480888
rect 169812 480848 170036 480876
rect 169812 480836 169818 480848
rect 170030 480836 170036 480848
rect 170088 480836 170094 480888
rect 173894 480836 173900 480888
rect 173952 480876 173958 480888
rect 174262 480876 174268 480888
rect 173952 480848 174268 480876
rect 173952 480836 173958 480848
rect 174262 480836 174268 480848
rect 174320 480836 174326 480888
rect 179414 480836 179420 480888
rect 179472 480876 179478 480888
rect 180058 480876 180064 480888
rect 179472 480848 180064 480876
rect 179472 480836 179478 480848
rect 180058 480836 180064 480848
rect 180116 480836 180122 480888
rect 182266 480836 182272 480888
rect 182324 480876 182330 480888
rect 183094 480876 183100 480888
rect 182324 480848 183100 480876
rect 182324 480836 182330 480848
rect 183094 480836 183100 480848
rect 183152 480836 183158 480888
rect 186314 480836 186320 480888
rect 186372 480876 186378 480888
rect 187142 480876 187148 480888
rect 186372 480848 187148 480876
rect 186372 480836 186378 480848
rect 187142 480836 187148 480848
rect 187200 480836 187206 480888
rect 205818 480836 205824 480888
rect 205876 480876 205882 480888
rect 206462 480876 206468 480888
rect 205876 480848 206468 480876
rect 205876 480836 205882 480848
rect 206462 480836 206468 480848
rect 206520 480836 206526 480888
rect 207198 480836 207204 480888
rect 207256 480876 207262 480888
rect 207566 480876 207572 480888
rect 207256 480848 207572 480876
rect 207256 480836 207262 480848
rect 207566 480836 207572 480848
rect 207624 480836 207630 480888
rect 209774 480836 209780 480888
rect 209832 480876 209838 480888
rect 209958 480876 209964 480888
rect 209832 480848 209964 480876
rect 209832 480836 209838 480848
rect 209958 480836 209964 480848
rect 210016 480836 210022 480888
rect 212534 480836 212540 480888
rect 212592 480876 212598 480888
rect 213454 480876 213460 480888
rect 212592 480848 213460 480876
rect 212592 480836 212598 480848
rect 213454 480836 213460 480848
rect 213512 480836 213518 480888
rect 248414 480836 248420 480888
rect 248472 480876 248478 480888
rect 249150 480876 249156 480888
rect 248472 480848 249156 480876
rect 248472 480836 248478 480848
rect 249150 480836 249156 480848
rect 249208 480836 249214 480888
rect 249886 480836 249892 480888
rect 249944 480876 249950 480888
rect 250070 480876 250076 480888
rect 249944 480848 250076 480876
rect 249944 480836 249950 480848
rect 250070 480836 250076 480848
rect 250128 480836 250134 480888
rect 251174 480836 251180 480888
rect 251232 480876 251238 480888
rect 251910 480876 251916 480888
rect 251232 480848 251916 480876
rect 251232 480836 251238 480848
rect 251910 480836 251916 480848
rect 251968 480836 251974 480888
rect 253934 480836 253940 480888
rect 253992 480876 253998 480888
rect 254118 480876 254124 480888
rect 253992 480848 254124 480876
rect 253992 480836 253998 480848
rect 254118 480836 254124 480848
rect 254176 480836 254182 480888
rect 262306 480836 262312 480888
rect 262364 480876 262370 480888
rect 262858 480876 262864 480888
rect 262364 480848 262864 480876
rect 262364 480836 262370 480848
rect 262858 480836 262864 480848
rect 262916 480836 262922 480888
rect 292574 480836 292580 480888
rect 292632 480876 292638 480888
rect 293310 480876 293316 480888
rect 292632 480848 293316 480876
rect 292632 480836 292638 480848
rect 293310 480836 293316 480848
rect 293368 480836 293374 480888
rect 293954 480836 293960 480888
rect 294012 480876 294018 480888
rect 294598 480876 294604 480888
rect 294012 480848 294604 480876
rect 294012 480836 294018 480848
rect 294598 480836 294604 480848
rect 294656 480836 294662 480888
rect 295518 480836 295524 480888
rect 295576 480876 295582 480888
rect 296254 480876 296260 480888
rect 295576 480848 296260 480876
rect 295576 480836 295582 480848
rect 296254 480836 296260 480848
rect 296312 480836 296318 480888
rect 70486 480768 70492 480820
rect 70544 480808 70550 480820
rect 71222 480808 71228 480820
rect 70544 480780 71228 480808
rect 70544 480768 70550 480780
rect 71222 480768 71228 480780
rect 71280 480768 71286 480820
rect 131206 480632 131212 480684
rect 131264 480672 131270 480684
rect 131574 480672 131580 480684
rect 131264 480644 131580 480672
rect 131264 480632 131270 480644
rect 131574 480632 131580 480644
rect 131632 480632 131638 480684
rect 171134 480292 171140 480344
rect 171192 480332 171198 480344
rect 171686 480332 171692 480344
rect 171192 480304 171692 480332
rect 171192 480292 171198 480304
rect 171686 480292 171692 480304
rect 171744 480292 171750 480344
rect 51718 480156 51724 480208
rect 51776 480196 51782 480208
rect 116118 480196 116124 480208
rect 51776 480168 116124 480196
rect 51776 480156 51782 480168
rect 116118 480156 116124 480168
rect 116176 480156 116182 480208
rect 292758 480156 292764 480208
rect 292816 480196 292822 480208
rect 368290 480196 368296 480208
rect 292816 480168 368296 480196
rect 292816 480156 292822 480168
rect 368290 480156 368296 480168
rect 368348 480156 368354 480208
rect 47394 480088 47400 480140
rect 47452 480128 47458 480140
rect 117590 480128 117596 480140
rect 47452 480100 117596 480128
rect 47452 480088 47458 480100
rect 117590 480088 117596 480100
rect 117648 480088 117654 480140
rect 281718 480088 281724 480140
rect 281776 480128 281782 480140
rect 359642 480128 359648 480140
rect 281776 480100 359648 480128
rect 281776 480088 281782 480100
rect 359642 480088 359648 480100
rect 359700 480088 359706 480140
rect 59630 480020 59636 480072
rect 59688 480060 59694 480072
rect 129918 480060 129924 480072
rect 59688 480032 129924 480060
rect 59688 480020 59694 480032
rect 129918 480020 129924 480032
rect 129976 480020 129982 480072
rect 297726 480020 297732 480072
rect 297784 480060 297790 480072
rect 376570 480060 376576 480072
rect 297784 480032 376576 480060
rect 297784 480020 297790 480032
rect 376570 480020 376576 480032
rect 376628 480020 376634 480072
rect 48958 479952 48964 480004
rect 49016 479992 49022 480004
rect 121546 479992 121552 480004
rect 49016 479964 121552 479992
rect 49016 479952 49022 479964
rect 121546 479952 121552 479964
rect 121604 479952 121610 480004
rect 278866 479952 278872 480004
rect 278924 479992 278930 480004
rect 364150 479992 364156 480004
rect 278924 479964 364156 479992
rect 278924 479952 278930 479964
rect 364150 479952 364156 479964
rect 364208 479952 364214 480004
rect 49142 479884 49148 479936
rect 49200 479924 49206 479936
rect 127710 479924 127716 479936
rect 49200 479896 127716 479924
rect 49200 479884 49206 479896
rect 127710 479884 127716 479896
rect 127768 479884 127774 479936
rect 275186 479884 275192 479936
rect 275244 479924 275250 479936
rect 370314 479924 370320 479936
rect 275244 479896 370320 479924
rect 275244 479884 275250 479896
rect 370314 479884 370320 479896
rect 370372 479884 370378 479936
rect 42518 479816 42524 479868
rect 42576 479856 42582 479868
rect 122926 479856 122932 479868
rect 42576 479828 122932 479856
rect 42576 479816 42582 479828
rect 122926 479816 122932 479828
rect 122984 479816 122990 479868
rect 260926 479816 260932 479868
rect 260984 479856 260990 479868
rect 368014 479856 368020 479868
rect 260984 479828 368020 479856
rect 260984 479816 260990 479828
rect 368014 479816 368020 479828
rect 368072 479816 368078 479868
rect 42426 479748 42432 479800
rect 42484 479788 42490 479800
rect 123294 479788 123300 479800
rect 42484 479760 123300 479788
rect 42484 479748 42490 479760
rect 123294 479748 123300 479760
rect 123352 479748 123358 479800
rect 265250 479748 265256 479800
rect 265308 479788 265314 479800
rect 373442 479788 373448 479800
rect 265308 479760 373448 479788
rect 265308 479748 265314 479760
rect 373442 479748 373448 479760
rect 373500 479748 373506 479800
rect 48866 479680 48872 479732
rect 48924 479720 48930 479732
rect 129734 479720 129740 479732
rect 48924 479692 129740 479720
rect 48924 479680 48930 479692
rect 129734 479680 129740 479692
rect 129792 479680 129798 479732
rect 254486 479680 254492 479732
rect 254544 479720 254550 479732
rect 366726 479720 366732 479732
rect 254544 479692 366732 479720
rect 254544 479680 254550 479692
rect 366726 479680 366732 479692
rect 366784 479680 366790 479732
rect 42334 479612 42340 479664
rect 42392 479652 42398 479664
rect 124582 479652 124588 479664
rect 42392 479624 124588 479652
rect 42392 479612 42398 479624
rect 124582 479612 124588 479624
rect 124640 479612 124646 479664
rect 253198 479612 253204 479664
rect 253256 479652 253262 479664
rect 374914 479652 374920 479664
rect 253256 479624 374920 479652
rect 253256 479612 253262 479624
rect 374914 479612 374920 479624
rect 374972 479612 374978 479664
rect 46106 479544 46112 479596
rect 46164 479584 46170 479596
rect 128998 479584 129004 479596
rect 46164 479556 129004 479584
rect 46164 479544 46170 479556
rect 128998 479544 129004 479556
rect 129056 479544 129062 479596
rect 158990 479544 158996 479596
rect 159048 479584 159054 479596
rect 207658 479584 207664 479596
rect 159048 479556 207664 479584
rect 159048 479544 159054 479556
rect 207658 479544 207664 479556
rect 207716 479544 207722 479596
rect 242986 479544 242992 479596
rect 243044 479584 243050 479596
rect 366542 479584 366548 479596
rect 243044 479556 366548 479584
rect 243044 479544 243050 479556
rect 366542 479544 366548 479556
rect 366600 479544 366606 479596
rect 62390 479476 62396 479528
rect 62448 479516 62454 479528
rect 199194 479516 199200 479528
rect 62448 479488 199200 479516
rect 62448 479476 62454 479488
rect 199194 479476 199200 479488
rect 199252 479476 199258 479528
rect 246482 479476 246488 479528
rect 246540 479516 246546 479528
rect 369302 479516 369308 479528
rect 246540 479488 369308 479516
rect 246540 479476 246546 479488
rect 369302 479476 369308 479488
rect 369360 479476 369366 479528
rect 54478 479408 54484 479460
rect 54536 479448 54542 479460
rect 117406 479448 117412 479460
rect 54536 479420 117412 479448
rect 54536 479408 54542 479420
rect 117406 479408 117412 479420
rect 117464 479408 117470 479460
rect 53282 479340 53288 479392
rect 53340 479380 53346 479392
rect 116210 479380 116216 479392
rect 53340 479352 116216 479380
rect 53340 479340 53346 479352
rect 116210 479340 116216 479352
rect 116268 479340 116274 479392
rect 53374 479272 53380 479324
rect 53432 479312 53438 479324
rect 116670 479312 116676 479324
rect 53432 479284 116676 479312
rect 53432 479272 53438 479284
rect 116670 479272 116676 479284
rect 116728 479272 116734 479324
rect 85574 479136 85580 479188
rect 85632 479176 85638 479188
rect 86310 479176 86316 479188
rect 85632 479148 86316 479176
rect 85632 479136 85638 479148
rect 86310 479136 86316 479148
rect 86368 479136 86374 479188
rect 169846 478728 169852 478780
rect 169904 478768 169910 478780
rect 170398 478768 170404 478780
rect 169904 478740 170404 478768
rect 169904 478728 169910 478740
rect 170398 478728 170404 478740
rect 170456 478728 170462 478780
rect 291470 478592 291476 478644
rect 291528 478632 291534 478644
rect 361390 478632 361396 478644
rect 291528 478604 361396 478632
rect 291528 478592 291534 478604
rect 361390 478592 361396 478604
rect 361448 478592 361454 478644
rect 288894 478524 288900 478576
rect 288952 478564 288958 478576
rect 361482 478564 361488 478576
rect 288952 478536 361488 478564
rect 288952 478524 288958 478536
rect 361482 478524 361488 478536
rect 361540 478524 361546 478576
rect 298462 478456 298468 478508
rect 298520 478496 298526 478508
rect 379238 478496 379244 478508
rect 298520 478468 379244 478496
rect 298520 478456 298526 478468
rect 379238 478456 379244 478468
rect 379296 478456 379302 478508
rect 244246 478400 253934 478428
rect 178126 478252 178132 478304
rect 178184 478292 178190 478304
rect 210694 478292 210700 478304
rect 178184 478264 210700 478292
rect 178184 478252 178190 478264
rect 210694 478252 210700 478264
rect 210752 478252 210758 478304
rect 238202 478252 238208 478304
rect 238260 478292 238266 478304
rect 244246 478292 244274 478400
rect 247402 478320 247408 478372
rect 247460 478360 247466 478372
rect 247460 478332 250760 478360
rect 247460 478320 247466 478332
rect 238260 478264 244274 478292
rect 238260 478252 238266 478264
rect 160186 478184 160192 478236
rect 160244 478224 160250 478236
rect 203518 478224 203524 478236
rect 160244 478196 203524 478224
rect 160244 478184 160250 478196
rect 203518 478184 203524 478196
rect 203576 478184 203582 478236
rect 249794 478184 249800 478236
rect 249852 478224 249858 478236
rect 250530 478224 250536 478236
rect 249852 478196 250536 478224
rect 249852 478184 249858 478196
rect 250530 478184 250536 478196
rect 250588 478184 250594 478236
rect 250732 478224 250760 478332
rect 253906 478292 253934 478400
rect 275646 478388 275652 478440
rect 275704 478428 275710 478440
rect 373718 478428 373724 478440
rect 275704 478400 373724 478428
rect 275704 478388 275710 478400
rect 373718 478388 373724 478400
rect 373776 478388 373782 478440
rect 260190 478320 260196 478372
rect 260248 478360 260254 478372
rect 370774 478360 370780 478372
rect 260248 478332 370780 478360
rect 260248 478320 260254 478332
rect 370774 478320 370780 478332
rect 370832 478320 370838 478372
rect 365070 478292 365076 478304
rect 253906 478264 365076 478292
rect 365070 478252 365076 478264
rect 365128 478252 365134 478304
rect 376018 478224 376024 478236
rect 250732 478196 376024 478224
rect 376018 478184 376024 478196
rect 376076 478184 376082 478236
rect 85666 478116 85672 478168
rect 85724 478156 85730 478168
rect 85850 478156 85856 478168
rect 85724 478128 85856 478156
rect 85724 478116 85730 478128
rect 85850 478116 85856 478128
rect 85908 478116 85914 478168
rect 146294 478116 146300 478168
rect 146352 478156 146358 478168
rect 218698 478156 218704 478168
rect 146352 478128 218704 478156
rect 146352 478116 146358 478128
rect 218698 478116 218704 478128
rect 218756 478116 218762 478168
rect 238754 478116 238760 478168
rect 238812 478156 238818 478168
rect 378870 478156 378876 478168
rect 238812 478128 378876 478156
rect 238812 478116 238818 478128
rect 378870 478116 378876 478128
rect 378928 478116 378934 478168
rect 273346 477844 273352 477896
rect 273404 477884 273410 477896
rect 273806 477884 273812 477896
rect 273404 477856 273812 477884
rect 273404 477844 273410 477856
rect 273806 477844 273812 477856
rect 273864 477844 273870 477896
rect 277394 477844 277400 477896
rect 277452 477884 277458 477896
rect 277854 477884 277860 477896
rect 277452 477856 277860 477884
rect 277452 477844 277458 477856
rect 277854 477844 277860 477856
rect 277912 477844 277918 477896
rect 78766 477640 78772 477692
rect 78824 477680 78830 477692
rect 79134 477680 79140 477692
rect 78824 477652 79140 477680
rect 78824 477640 78830 477652
rect 79134 477640 79140 477652
rect 79192 477640 79198 477692
rect 59722 477436 59728 477488
rect 59780 477476 59786 477488
rect 133874 477476 133880 477488
rect 59780 477448 133880 477476
rect 59780 477436 59786 477448
rect 133874 477436 133880 477448
rect 133932 477436 133938 477488
rect 46842 477368 46848 477420
rect 46900 477408 46906 477420
rect 122834 477408 122840 477420
rect 46900 477380 122840 477408
rect 46900 477368 46906 477380
rect 122834 477368 122840 477380
rect 122892 477368 122898 477420
rect 207106 477368 207112 477420
rect 207164 477408 207170 477420
rect 207750 477408 207756 477420
rect 207164 477380 207756 477408
rect 207164 477368 207170 477380
rect 207750 477368 207756 477380
rect 207808 477368 207814 477420
rect 291286 477368 291292 477420
rect 291344 477408 291350 477420
rect 365530 477408 365536 477420
rect 291344 477380 365536 477408
rect 291344 477368 291350 477380
rect 365530 477368 365536 477380
rect 365588 477368 365594 477420
rect 57330 477300 57336 477352
rect 57388 477340 57394 477352
rect 135990 477340 135996 477352
rect 57388 477312 135996 477340
rect 57388 477300 57394 477312
rect 135990 477300 135996 477312
rect 136048 477300 136054 477352
rect 276566 477300 276572 477352
rect 276624 477340 276630 477352
rect 358722 477340 358728 477352
rect 276624 477312 358728 477340
rect 276624 477300 276630 477312
rect 358722 477300 358728 477312
rect 358780 477300 358786 477352
rect 55766 477232 55772 477284
rect 55824 477272 55830 477284
rect 134702 477272 134708 477284
rect 55824 477244 134708 477272
rect 55824 477232 55830 477244
rect 134702 477232 134708 477244
rect 134760 477232 134766 477284
rect 274726 477232 274732 477284
rect 274784 477272 274790 477284
rect 365438 477272 365444 477284
rect 274784 477244 365444 477272
rect 274784 477232 274790 477244
rect 365438 477232 365444 477244
rect 365496 477232 365502 477284
rect 50154 477164 50160 477216
rect 50212 477204 50218 477216
rect 131298 477204 131304 477216
rect 50212 477176 131304 477204
rect 50212 477164 50218 477176
rect 131298 477164 131304 477176
rect 131356 477164 131362 477216
rect 264238 477164 264244 477216
rect 264296 477204 264302 477216
rect 362586 477204 362592 477216
rect 264296 477176 362592 477204
rect 264296 477164 264302 477176
rect 362586 477164 362592 477176
rect 362644 477164 362650 477216
rect 47854 477096 47860 477148
rect 47912 477136 47918 477148
rect 129826 477136 129832 477148
rect 47912 477108 129832 477136
rect 47912 477096 47918 477108
rect 129826 477096 129832 477108
rect 129884 477096 129890 477148
rect 263594 477096 263600 477148
rect 263652 477136 263658 477148
rect 363966 477136 363972 477148
rect 263652 477108 363972 477136
rect 263652 477096 263658 477108
rect 363966 477096 363972 477108
rect 364024 477096 364030 477148
rect 48774 477028 48780 477080
rect 48832 477068 48838 477080
rect 133414 477068 133420 477080
rect 48832 477040 133420 477068
rect 48832 477028 48838 477040
rect 133414 477028 133420 477040
rect 133472 477028 133478 477080
rect 263686 477028 263692 477080
rect 263744 477068 263750 477080
rect 365346 477068 365352 477080
rect 263744 477040 365352 477068
rect 263744 477028 263750 477040
rect 365346 477028 365352 477040
rect 365404 477028 365410 477080
rect 46198 476960 46204 477012
rect 46256 477000 46262 477012
rect 132586 477000 132592 477012
rect 46256 476972 132592 477000
rect 46256 476960 46262 476972
rect 132586 476960 132592 476972
rect 132644 476960 132650 477012
rect 204530 476960 204536 477012
rect 204588 477000 204594 477012
rect 217318 477000 217324 477012
rect 204588 476972 217324 477000
rect 204588 476960 204594 476972
rect 217318 476960 217324 476972
rect 217376 476960 217382 477012
rect 259730 476960 259736 477012
rect 259788 477000 259794 477012
rect 363874 477000 363880 477012
rect 259788 476972 363880 477000
rect 259788 476960 259794 476972
rect 363874 476960 363880 476972
rect 363932 476960 363938 477012
rect 43990 476892 43996 476944
rect 44048 476932 44054 476944
rect 132494 476932 132500 476944
rect 44048 476904 132500 476932
rect 44048 476892 44054 476904
rect 132494 476892 132500 476904
rect 132552 476892 132558 476944
rect 188062 476892 188068 476944
rect 188120 476932 188126 476944
rect 207750 476932 207756 476944
rect 188120 476904 207756 476932
rect 188120 476892 188126 476904
rect 207750 476892 207756 476904
rect 207808 476892 207814 476944
rect 258534 476892 258540 476944
rect 258592 476932 258598 476944
rect 368106 476932 368112 476944
rect 258592 476904 368112 476932
rect 258592 476892 258598 476904
rect 368106 476892 368112 476904
rect 368164 476892 368170 476944
rect 45002 476824 45008 476876
rect 45060 476864 45066 476876
rect 133966 476864 133972 476876
rect 45060 476836 133972 476864
rect 45060 476824 45066 476836
rect 133966 476824 133972 476836
rect 134024 476824 134030 476876
rect 185762 476824 185768 476876
rect 185820 476864 185826 476876
rect 213270 476864 213276 476876
rect 185820 476836 213276 476864
rect 185820 476824 185826 476836
rect 213270 476824 213276 476836
rect 213328 476824 213334 476876
rect 246114 476824 246120 476876
rect 246172 476864 246178 476876
rect 362402 476864 362408 476876
rect 246172 476836 362408 476864
rect 246172 476824 246178 476836
rect 362402 476824 362408 476836
rect 362460 476824 362466 476876
rect 44726 476756 44732 476808
rect 44784 476796 44790 476808
rect 143718 476796 143724 476808
rect 44784 476768 143724 476796
rect 44784 476756 44790 476768
rect 143718 476756 143724 476768
rect 143776 476756 143782 476808
rect 164602 476756 164608 476808
rect 164660 476796 164666 476808
rect 211890 476796 211896 476808
rect 164660 476768 211896 476796
rect 164660 476756 164666 476768
rect 211890 476756 211896 476768
rect 211948 476756 211954 476808
rect 244458 476756 244464 476808
rect 244516 476796 244522 476808
rect 373258 476796 373264 476808
rect 244516 476768 373264 476796
rect 244516 476756 244522 476768
rect 373258 476756 373264 476768
rect 373316 476756 373322 476808
rect 57146 476688 57152 476740
rect 57204 476728 57210 476740
rect 131206 476728 131212 476740
rect 57204 476700 131212 476728
rect 57204 476688 57210 476700
rect 131206 476688 131212 476700
rect 131264 476688 131270 476740
rect 58434 476620 58440 476672
rect 58492 476660 58498 476672
rect 131114 476660 131120 476672
rect 58492 476632 131120 476660
rect 58492 476620 58498 476632
rect 131114 476620 131120 476632
rect 131172 476620 131178 476672
rect 58526 476552 58532 476604
rect 58584 476592 58590 476604
rect 128446 476592 128452 476604
rect 58584 476564 128452 476592
rect 58584 476552 58590 476564
rect 128446 476552 128452 476564
rect 128504 476552 128510 476604
rect 175274 476416 175280 476468
rect 175332 476456 175338 476468
rect 176102 476456 176108 476468
rect 175332 476428 176108 476456
rect 175332 476416 175338 476428
rect 176102 476416 176108 476428
rect 176160 476416 176166 476468
rect 278774 475804 278780 475856
rect 278832 475844 278838 475856
rect 357066 475844 357072 475856
rect 278832 475816 357072 475844
rect 278832 475804 278838 475816
rect 357066 475804 357072 475816
rect 357124 475804 357130 475856
rect 270862 475736 270868 475788
rect 270920 475776 270926 475788
rect 364242 475776 364248 475788
rect 270920 475748 364248 475776
rect 270920 475736 270926 475748
rect 364242 475736 364248 475748
rect 364300 475736 364306 475788
rect 274634 475668 274640 475720
rect 274692 475708 274698 475720
rect 368382 475708 368388 475720
rect 274692 475680 368388 475708
rect 274692 475668 274698 475680
rect 368382 475668 368388 475680
rect 368440 475668 368446 475720
rect 187786 475600 187792 475652
rect 187844 475640 187850 475652
rect 200942 475640 200948 475652
rect 187844 475612 200948 475640
rect 187844 475600 187850 475612
rect 200942 475600 200948 475612
rect 201000 475600 201006 475652
rect 259454 475600 259460 475652
rect 259512 475640 259518 475652
rect 372246 475640 372252 475652
rect 259512 475612 372252 475640
rect 259512 475600 259518 475612
rect 372246 475600 372252 475612
rect 372304 475600 372310 475652
rect 179598 475532 179604 475584
rect 179656 475572 179662 475584
rect 219066 475572 219072 475584
rect 179656 475544 219072 475572
rect 179656 475532 179662 475544
rect 219066 475532 219072 475544
rect 219124 475532 219130 475584
rect 236454 475532 236460 475584
rect 236512 475572 236518 475584
rect 362310 475572 362316 475584
rect 236512 475544 362316 475572
rect 236512 475532 236518 475544
rect 362310 475532 362316 475544
rect 362368 475532 362374 475584
rect 162946 475464 162952 475516
rect 163004 475504 163010 475516
rect 206370 475504 206376 475516
rect 163004 475476 206376 475504
rect 163004 475464 163010 475476
rect 206370 475464 206376 475476
rect 206428 475464 206434 475516
rect 232406 475464 232412 475516
rect 232464 475504 232470 475516
rect 367738 475504 367744 475516
rect 232464 475476 367744 475504
rect 232464 475464 232470 475476
rect 367738 475464 367744 475476
rect 367796 475464 367802 475516
rect 168650 475396 168656 475448
rect 168708 475436 168714 475448
rect 213178 475436 213184 475448
rect 168708 475408 213184 475436
rect 168708 475396 168714 475408
rect 213178 475396 213184 475408
rect 213236 475396 213242 475448
rect 237466 475396 237472 475448
rect 237524 475436 237530 475448
rect 376110 475436 376116 475448
rect 237524 475408 376116 475436
rect 237524 475396 237530 475408
rect 376110 475396 376116 475408
rect 376168 475396 376174 475448
rect 61010 475328 61016 475380
rect 61068 475368 61074 475380
rect 199562 475368 199568 475380
rect 61068 475340 199568 475368
rect 61068 475328 61074 475340
rect 199562 475328 199568 475340
rect 199620 475328 199626 475380
rect 206094 475328 206100 475380
rect 206152 475368 206158 475380
rect 217686 475368 217692 475380
rect 206152 475340 217692 475368
rect 206152 475328 206158 475340
rect 217686 475328 217692 475340
rect 217744 475328 217750 475380
rect 229186 475328 229192 475380
rect 229244 475368 229250 475380
rect 369118 475368 369124 475380
rect 229244 475340 369124 475368
rect 229244 475328 229250 475340
rect 369118 475328 369124 475340
rect 369176 475328 369182 475380
rect 45370 474512 45376 474564
rect 45428 474552 45434 474564
rect 73890 474552 73896 474564
rect 45428 474524 73896 474552
rect 45428 474512 45434 474524
rect 73890 474512 73896 474524
rect 73948 474512 73954 474564
rect 54754 474444 54760 474496
rect 54812 474484 54818 474496
rect 101582 474484 101588 474496
rect 54812 474456 101588 474484
rect 54812 474444 54818 474456
rect 101582 474444 101588 474456
rect 101640 474444 101646 474496
rect 289906 474444 289912 474496
rect 289964 474484 289970 474496
rect 367002 474484 367008 474496
rect 289964 474456 367008 474484
rect 289964 474444 289970 474456
rect 367002 474444 367008 474456
rect 367060 474444 367066 474496
rect 53190 474376 53196 474428
rect 53248 474416 53254 474428
rect 99926 474416 99932 474428
rect 53248 474388 99932 474416
rect 53248 474376 53254 474388
rect 99926 474376 99932 474388
rect 99984 474376 99990 474428
rect 290182 474376 290188 474428
rect 290240 474416 290246 474428
rect 374454 474416 374460 474428
rect 290240 474388 374460 474416
rect 290240 474376 290246 474388
rect 374454 474376 374460 474388
rect 374512 474376 374518 474428
rect 57422 474308 57428 474360
rect 57480 474348 57486 474360
rect 103698 474348 103704 474360
rect 57480 474320 103704 474348
rect 57480 474308 57486 474320
rect 103698 474308 103704 474320
rect 103756 474308 103762 474360
rect 178034 474308 178040 474360
rect 178092 474348 178098 474360
rect 202138 474348 202144 474360
rect 178092 474320 202144 474348
rect 178092 474308 178098 474320
rect 202138 474308 202144 474320
rect 202196 474308 202202 474360
rect 273438 474308 273444 474360
rect 273496 474348 273502 474360
rect 360746 474348 360752 474360
rect 273496 474320 360752 474348
rect 273496 474308 273502 474320
rect 360746 474308 360752 474320
rect 360804 474308 360810 474360
rect 50338 474240 50344 474292
rect 50396 474280 50402 474292
rect 98638 474280 98644 474292
rect 50396 474252 98644 474280
rect 50396 474240 50402 474252
rect 98638 474240 98644 474252
rect 98696 474240 98702 474292
rect 172054 474240 172060 474292
rect 172112 474280 172118 474292
rect 210510 474280 210516 474292
rect 172112 474252 210516 474280
rect 172112 474240 172118 474252
rect 210510 474240 210516 474252
rect 210568 474240 210574 474292
rect 257614 474240 257620 474292
rect 257672 474280 257678 474292
rect 366818 474280 366824 474292
rect 257672 474252 366824 474280
rect 257672 474240 257678 474252
rect 366818 474240 366824 474252
rect 366876 474240 366882 474292
rect 51534 474172 51540 474224
rect 51592 474212 51598 474224
rect 99466 474212 99472 474224
rect 51592 474184 99472 474212
rect 51592 474172 51598 474184
rect 99466 474172 99472 474184
rect 99524 474172 99530 474224
rect 158714 474172 158720 474224
rect 158772 474212 158778 474224
rect 209038 474212 209044 474224
rect 158772 474184 209044 474212
rect 158772 474172 158778 474184
rect 209038 474172 209044 474184
rect 209096 474172 209102 474224
rect 262398 474172 262404 474224
rect 262456 474212 262462 474224
rect 373534 474212 373540 474224
rect 262456 474184 373540 474212
rect 262456 474172 262462 474184
rect 373534 474172 373540 474184
rect 373592 474172 373598 474224
rect 57698 474104 57704 474156
rect 57756 474144 57762 474156
rect 113542 474144 113548 474156
rect 57756 474116 113548 474144
rect 57756 474104 57762 474116
rect 113542 474104 113548 474116
rect 113600 474104 113606 474156
rect 153194 474104 153200 474156
rect 153252 474144 153258 474156
rect 218790 474144 218796 474156
rect 153252 474116 218796 474144
rect 153252 474104 153258 474116
rect 218790 474104 218796 474116
rect 218848 474104 218854 474156
rect 244366 474104 244372 474156
rect 244424 474144 244430 474156
rect 360930 474144 360936 474156
rect 244424 474116 360936 474144
rect 244424 474104 244430 474116
rect 360930 474104 360936 474116
rect 360988 474104 360994 474156
rect 45278 474036 45284 474088
rect 45336 474076 45342 474088
rect 106366 474076 106372 474088
rect 45336 474048 106372 474076
rect 45336 474036 45342 474048
rect 106366 474036 106372 474048
rect 106424 474036 106430 474088
rect 139486 474036 139492 474088
rect 139544 474076 139550 474088
rect 207290 474076 207296 474088
rect 139544 474048 207296 474076
rect 139544 474036 139550 474048
rect 207290 474036 207296 474048
rect 207348 474036 207354 474088
rect 240134 474036 240140 474088
rect 240192 474076 240198 474088
rect 369394 474076 369400 474088
rect 240192 474048 369400 474076
rect 240192 474036 240198 474048
rect 369394 474036 369400 474048
rect 369452 474036 369458 474088
rect 59354 473968 59360 474020
rect 59412 474008 59418 474020
rect 180150 474008 180156 474020
rect 59412 473980 180156 474008
rect 59412 473968 59418 473980
rect 180150 473968 180156 473980
rect 180208 473968 180214 474020
rect 186406 473968 186412 474020
rect 186464 474008 186470 474020
rect 212074 474008 212080 474020
rect 186464 473980 212080 474008
rect 186464 473968 186470 473980
rect 212074 473968 212080 473980
rect 212132 473968 212138 474020
rect 240778 473968 240784 474020
rect 240836 474008 240842 474020
rect 374638 474008 374644 474020
rect 240836 473980 374644 474008
rect 240836 473968 240842 473980
rect 374638 473968 374644 473980
rect 374696 473968 374702 474020
rect 291194 473152 291200 473204
rect 291252 473192 291258 473204
rect 357158 473192 357164 473204
rect 291252 473164 357164 473192
rect 291252 473152 291258 473164
rect 357158 473152 357164 473164
rect 357216 473152 357222 473204
rect 280154 473084 280160 473136
rect 280212 473124 280218 473136
rect 366266 473124 366272 473136
rect 280212 473096 366272 473124
rect 280212 473084 280218 473096
rect 366266 473084 366272 473096
rect 366324 473084 366330 473136
rect 273346 473016 273352 473068
rect 273404 473056 273410 473068
rect 362862 473056 362868 473068
rect 273404 473028 362868 473056
rect 273404 473016 273410 473028
rect 362862 473016 362868 473028
rect 362920 473016 362926 473068
rect 262306 472948 262312 473000
rect 262364 472988 262370 473000
rect 372338 472988 372344 473000
rect 262364 472960 372344 472988
rect 262364 472948 262370 472960
rect 372338 472948 372344 472960
rect 372396 472948 372402 473000
rect 258166 472880 258172 472932
rect 258224 472920 258230 472932
rect 370866 472920 370872 472932
rect 258224 472892 370872 472920
rect 258224 472880 258230 472892
rect 370866 472880 370872 472892
rect 370924 472880 370930 472932
rect 58710 472812 58716 472864
rect 58768 472852 58774 472864
rect 110598 472852 110604 472864
rect 58768 472824 110604 472852
rect 58768 472812 58774 472824
rect 110598 472812 110604 472824
rect 110656 472812 110662 472864
rect 241606 472812 241612 472864
rect 241664 472852 241670 472864
rect 376202 472852 376208 472864
rect 241664 472824 376208 472852
rect 241664 472812 241670 472824
rect 376202 472812 376208 472824
rect 376260 472812 376266 472864
rect 45186 472744 45192 472796
rect 45244 472784 45250 472796
rect 105630 472784 105636 472796
rect 45244 472756 105636 472784
rect 45244 472744 45250 472756
rect 105630 472744 105636 472756
rect 105688 472744 105694 472796
rect 226334 472744 226340 472796
rect 226392 472784 226398 472796
rect 364978 472784 364984 472796
rect 226392 472756 364984 472784
rect 226392 472744 226398 472756
rect 364978 472744 364984 472756
rect 365036 472744 365042 472796
rect 45094 472676 45100 472728
rect 45152 472716 45158 472728
rect 104986 472716 104992 472728
rect 45152 472688 104992 472716
rect 45152 472676 45158 472688
rect 104986 472676 104992 472688
rect 105044 472676 105050 472728
rect 175366 472676 175372 472728
rect 175424 472716 175430 472728
rect 210786 472716 210792 472728
rect 175424 472688 210792 472716
rect 175424 472676 175430 472688
rect 210786 472676 210792 472688
rect 210844 472676 210850 472728
rect 237374 472676 237380 472728
rect 237432 472716 237438 472728
rect 378962 472716 378968 472728
rect 237432 472688 378968 472716
rect 237432 472676 237438 472688
rect 378962 472676 378968 472688
rect 379020 472676 379026 472728
rect 43438 472608 43444 472660
rect 43496 472648 43502 472660
rect 103606 472648 103612 472660
rect 43496 472620 103612 472648
rect 43496 472608 43502 472620
rect 103606 472608 103612 472620
rect 103664 472608 103670 472660
rect 179506 472608 179512 472660
rect 179564 472648 179570 472660
rect 216214 472648 216220 472660
rect 179564 472620 216220 472648
rect 179564 472608 179570 472620
rect 216214 472608 216220 472620
rect 216272 472608 216278 472660
rect 227254 472608 227260 472660
rect 227312 472648 227318 472660
rect 371970 472648 371976 472660
rect 227312 472620 371976 472648
rect 227312 472608 227318 472620
rect 371970 472608 371976 472620
rect 372028 472608 372034 472660
rect 50890 471928 50896 471980
rect 50948 471968 50954 471980
rect 81894 471968 81900 471980
rect 50948 471940 81900 471968
rect 50948 471928 50954 471940
rect 81894 471928 81900 471940
rect 81952 471928 81958 471980
rect 185026 471928 185032 471980
rect 185084 471968 185090 471980
rect 206554 471968 206560 471980
rect 185084 471940 206560 471968
rect 185084 471928 185090 471940
rect 206554 471928 206560 471940
rect 206612 471928 206618 471980
rect 295886 471928 295892 471980
rect 295944 471968 295950 471980
rect 369762 471968 369768 471980
rect 295944 471940 369768 471968
rect 295944 471928 295950 471940
rect 369762 471928 369768 471940
rect 369820 471928 369826 471980
rect 53558 471860 53564 471912
rect 53616 471900 53622 471912
rect 84470 471900 84476 471912
rect 53616 471872 84476 471900
rect 53616 471860 53622 471872
rect 84470 471860 84476 471872
rect 84528 471860 84534 471912
rect 189718 471860 189724 471912
rect 189776 471900 189782 471912
rect 215018 471900 215024 471912
rect 189776 471872 215024 471900
rect 189776 471860 189782 471872
rect 215018 471860 215024 471872
rect 215076 471860 215082 471912
rect 295518 471860 295524 471912
rect 295576 471900 295582 471912
rect 370222 471900 370228 471912
rect 295576 471872 370228 471900
rect 295576 471860 295582 471872
rect 370222 471860 370228 471872
rect 370280 471860 370286 471912
rect 50798 471792 50804 471844
rect 50856 471832 50862 471844
rect 82814 471832 82820 471844
rect 50856 471804 82820 471832
rect 50856 471792 50862 471804
rect 82814 471792 82820 471804
rect 82872 471792 82878 471844
rect 191006 471792 191012 471844
rect 191064 471832 191070 471844
rect 217410 471832 217416 471844
rect 191064 471804 217416 471832
rect 191064 471792 191070 471804
rect 217410 471792 217416 471804
rect 217468 471792 217474 471844
rect 295426 471792 295432 471844
rect 295484 471832 295490 471844
rect 371234 471832 371240 471844
rect 295484 471804 371240 471832
rect 295484 471792 295490 471804
rect 371234 471792 371240 471804
rect 371292 471792 371298 471844
rect 51442 471724 51448 471776
rect 51500 471764 51506 471776
rect 84286 471764 84292 471776
rect 51500 471736 84292 471764
rect 51500 471724 51506 471736
rect 84286 471724 84292 471736
rect 84344 471724 84350 471776
rect 181438 471724 181444 471776
rect 181496 471764 181502 471776
rect 209314 471764 209320 471776
rect 181496 471736 209320 471764
rect 181496 471724 181502 471736
rect 209314 471724 209320 471736
rect 209372 471724 209378 471776
rect 288434 471724 288440 471776
rect 288492 471764 288498 471776
rect 364886 471764 364892 471776
rect 288492 471736 364892 471764
rect 288492 471724 288498 471736
rect 364886 471724 364892 471736
rect 364944 471724 364950 471776
rect 53650 471656 53656 471708
rect 53708 471696 53714 471708
rect 85758 471696 85764 471708
rect 53708 471668 85764 471696
rect 53708 471656 53714 471668
rect 85758 471656 85764 471668
rect 85816 471656 85822 471708
rect 182726 471656 182732 471708
rect 182784 471696 182790 471708
rect 210878 471696 210884 471708
rect 182784 471668 210884 471696
rect 182784 471656 182790 471668
rect 210878 471656 210884 471668
rect 210936 471656 210942 471708
rect 296714 471656 296720 471708
rect 296772 471696 296778 471708
rect 373810 471696 373816 471708
rect 296772 471668 373816 471696
rect 296772 471656 296778 471668
rect 373810 471656 373816 471668
rect 373868 471656 373874 471708
rect 50706 471588 50712 471640
rect 50764 471628 50770 471640
rect 82906 471628 82912 471640
rect 50764 471600 82912 471628
rect 50764 471588 50770 471600
rect 82906 471588 82912 471600
rect 82964 471588 82970 471640
rect 182266 471588 182272 471640
rect 182324 471628 182330 471640
rect 216306 471628 216312 471640
rect 182324 471600 216312 471628
rect 182324 471588 182330 471600
rect 216306 471588 216312 471600
rect 216364 471588 216370 471640
rect 298094 471588 298100 471640
rect 298152 471628 298158 471640
rect 375374 471628 375380 471640
rect 298152 471600 375380 471628
rect 298152 471588 298158 471600
rect 375374 471588 375380 471600
rect 375432 471588 375438 471640
rect 49418 471520 49424 471572
rect 49476 471560 49482 471572
rect 83182 471560 83188 471572
rect 49476 471532 83188 471560
rect 49476 471520 49482 471532
rect 83182 471520 83188 471532
rect 83240 471520 83246 471572
rect 161658 471520 161664 471572
rect 161716 471560 161722 471572
rect 210602 471560 210608 471572
rect 161716 471532 210608 471560
rect 161716 471520 161722 471532
rect 210602 471520 210608 471532
rect 210660 471520 210666 471572
rect 295334 471520 295340 471572
rect 295392 471560 295398 471572
rect 377122 471560 377128 471572
rect 295392 471532 377128 471560
rect 295392 471520 295398 471532
rect 377122 471520 377128 471532
rect 377180 471520 377186 471572
rect 58894 471452 58900 471504
rect 58952 471492 58958 471504
rect 95510 471492 95516 471504
rect 58952 471464 95516 471492
rect 58952 471452 58958 471464
rect 95510 471452 95516 471464
rect 95568 471452 95574 471504
rect 140958 471452 140964 471504
rect 141016 471492 141022 471504
rect 200390 471492 200396 471504
rect 141016 471464 200396 471492
rect 141016 471452 141022 471464
rect 200390 471452 200396 471464
rect 200448 471452 200454 471504
rect 286134 471452 286140 471504
rect 286192 471492 286198 471504
rect 377950 471492 377956 471504
rect 286192 471464 377956 471492
rect 286192 471452 286198 471464
rect 377950 471452 377956 471464
rect 378008 471452 378014 471504
rect 53098 471384 53104 471436
rect 53156 471424 53162 471436
rect 100754 471424 100760 471436
rect 53156 471396 100760 471424
rect 53156 471384 53162 471396
rect 100754 471384 100760 471396
rect 100812 471384 100818 471436
rect 140866 471384 140872 471436
rect 140924 471424 140930 471436
rect 195238 471424 195244 471436
rect 140924 471396 195244 471424
rect 140924 471384 140930 471396
rect 195238 471384 195244 471396
rect 195296 471384 195302 471436
rect 195330 471384 195336 471436
rect 195388 471424 195394 471436
rect 200482 471424 200488 471436
rect 195388 471396 200488 471424
rect 195388 471384 195394 471396
rect 200482 471384 200488 471396
rect 200540 471384 200546 471436
rect 287146 471384 287152 471436
rect 287204 471424 287210 471436
rect 379330 471424 379336 471436
rect 287204 471396 379336 471424
rect 287204 471384 287210 471396
rect 379330 471384 379336 471396
rect 379388 471384 379394 471436
rect 57514 471316 57520 471368
rect 57572 471356 57578 471368
rect 114738 471356 114744 471368
rect 57572 471328 114744 471356
rect 57572 471316 57578 471328
rect 114738 471316 114744 471328
rect 114796 471316 114802 471368
rect 124214 471316 124220 471368
rect 124272 471356 124278 471368
rect 196894 471356 196900 471368
rect 124272 471328 196900 471356
rect 124272 471316 124278 471328
rect 196894 471316 196900 471328
rect 196952 471316 196958 471368
rect 255406 471316 255412 471368
rect 255464 471356 255470 471368
rect 358446 471356 358452 471368
rect 255464 471328 358452 471356
rect 255464 471316 255470 471328
rect 358446 471316 358452 471328
rect 358504 471316 358510 471368
rect 53006 471248 53012 471300
rect 53064 471288 53070 471300
rect 100846 471288 100852 471300
rect 53064 471260 100852 471288
rect 53064 471248 53070 471260
rect 100846 471248 100852 471260
rect 100904 471248 100910 471300
rect 108206 471248 108212 471300
rect 108264 471288 108270 471300
rect 202874 471288 202880 471300
rect 108264 471260 202880 471288
rect 108264 471248 108270 471260
rect 202874 471248 202880 471260
rect 202932 471248 202938 471300
rect 251358 471248 251364 471300
rect 251416 471288 251422 471300
rect 366634 471288 366640 471300
rect 251416 471260 366640 471288
rect 251416 471248 251422 471260
rect 366634 471248 366640 471260
rect 366692 471248 366698 471300
rect 44910 471180 44916 471232
rect 44968 471220 44974 471232
rect 65058 471220 65064 471232
rect 44968 471192 65064 471220
rect 44968 471180 44974 471192
rect 65058 471180 65064 471192
rect 65116 471180 65122 471232
rect 182358 471180 182364 471232
rect 182416 471220 182422 471232
rect 203702 471220 203708 471232
rect 182416 471192 203708 471220
rect 182416 471180 182422 471192
rect 203702 471180 203708 471192
rect 203760 471180 203766 471232
rect 287514 471180 287520 471232
rect 287572 471220 287578 471232
rect 359550 471220 359556 471232
rect 287572 471192 359556 471220
rect 287572 471180 287578 471192
rect 359550 471180 359556 471192
rect 359608 471180 359614 471232
rect 44818 471112 44824 471164
rect 44876 471152 44882 471164
rect 64874 471152 64880 471164
rect 44876 471124 64880 471152
rect 44876 471112 44882 471124
rect 64874 471112 64880 471124
rect 64932 471112 64938 471164
rect 185578 471112 185584 471164
rect 185636 471152 185642 471164
rect 205910 471152 205916 471164
rect 185636 471124 205916 471152
rect 185636 471112 185642 471124
rect 205910 471112 205916 471124
rect 205968 471112 205974 471164
rect 299474 471112 299480 471164
rect 299532 471152 299538 471164
rect 364794 471152 364800 471164
rect 299532 471124 364800 471152
rect 299532 471112 299538 471124
rect 364794 471112 364800 471124
rect 364852 471112 364858 471164
rect 47762 471044 47768 471096
rect 47820 471084 47826 471096
rect 64966 471084 64972 471096
rect 47820 471056 64972 471084
rect 47820 471044 47826 471056
rect 64966 471044 64972 471056
rect 65024 471044 65030 471096
rect 195238 471044 195244 471096
rect 195296 471084 195302 471096
rect 201862 471084 201868 471096
rect 195296 471056 201868 471084
rect 195296 471044 195302 471056
rect 201862 471044 201868 471056
rect 201920 471044 201926 471096
rect 193858 470976 193864 471028
rect 193916 471016 193922 471028
rect 195330 471016 195336 471028
rect 193916 470988 195336 471016
rect 193916 470976 193922 470988
rect 195330 470976 195336 470988
rect 195388 470976 195394 471028
rect 289814 470500 289820 470552
rect 289872 470540 289878 470552
rect 360654 470540 360660 470552
rect 289872 470512 360660 470540
rect 289872 470500 289878 470512
rect 360654 470500 360660 470512
rect 360712 470500 360718 470552
rect 283098 470432 283104 470484
rect 283156 470472 283162 470484
rect 358078 470472 358084 470484
rect 283156 470444 358084 470472
rect 283156 470432 283162 470444
rect 358078 470432 358084 470444
rect 358136 470432 358142 470484
rect 282914 470364 282920 470416
rect 282972 470404 282978 470416
rect 359918 470404 359924 470416
rect 282972 470376 359924 470404
rect 282972 470364 282978 470376
rect 359918 470364 359924 470376
rect 359976 470364 359982 470416
rect 283006 470296 283012 470348
rect 283064 470336 283070 470348
rect 360010 470336 360016 470348
rect 283064 470308 360016 470336
rect 283064 470296 283070 470308
rect 360010 470296 360016 470308
rect 360068 470296 360074 470348
rect 287054 470228 287060 470280
rect 287112 470268 287118 470280
rect 367554 470268 367560 470280
rect 287112 470240 367560 470268
rect 287112 470228 287118 470240
rect 367554 470228 367560 470240
rect 367612 470228 367618 470280
rect 285766 470160 285772 470212
rect 285824 470200 285830 470212
rect 373902 470200 373908 470212
rect 285824 470172 373908 470200
rect 285824 470160 285830 470172
rect 373902 470160 373908 470172
rect 373960 470160 373966 470212
rect 281534 470092 281540 470144
rect 281592 470132 281598 470144
rect 371142 470132 371148 470144
rect 281592 470104 371148 470132
rect 281592 470092 281598 470104
rect 371142 470092 371148 470104
rect 371200 470092 371206 470144
rect 270494 470024 270500 470076
rect 270552 470064 270558 470076
rect 362770 470064 362776 470076
rect 270552 470036 362776 470064
rect 270552 470024 270558 470036
rect 362770 470024 362776 470036
rect 362828 470024 362834 470076
rect 284386 469956 284392 470008
rect 284444 469996 284450 470008
rect 377490 469996 377496 470008
rect 284444 469968 377496 469996
rect 284444 469956 284450 469968
rect 377490 469956 377496 469968
rect 377548 469956 377554 470008
rect 172606 469888 172612 469940
rect 172664 469928 172670 469940
rect 205082 469928 205088 469940
rect 172664 469900 205088 469928
rect 172664 469888 172670 469900
rect 205082 469888 205088 469900
rect 205140 469888 205146 469940
rect 284294 469888 284300 469940
rect 284352 469928 284358 469940
rect 377582 469928 377588 469940
rect 284352 469900 377588 469928
rect 284352 469888 284358 469900
rect 377582 469888 377588 469900
rect 377640 469888 377646 469940
rect 57606 469820 57612 469872
rect 57664 469860 57670 469872
rect 111978 469860 111984 469872
rect 57664 469832 111984 469860
rect 57664 469820 57670 469832
rect 111978 469820 111984 469832
rect 112036 469820 112042 469872
rect 160094 469820 160100 469872
rect 160152 469860 160158 469872
rect 202322 469860 202328 469872
rect 160152 469832 202328 469860
rect 160152 469820 160158 469832
rect 202322 469820 202328 469832
rect 202380 469820 202386 469872
rect 281626 469820 281632 469872
rect 281684 469860 281690 469872
rect 379882 469860 379888 469872
rect 281684 469832 379888 469860
rect 281684 469820 281690 469832
rect 379882 469820 379888 469832
rect 379940 469820 379946 469872
rect 51350 469140 51356 469192
rect 51408 469180 51414 469192
rect 68278 469180 68284 469192
rect 51408 469152 68284 469180
rect 51408 469140 51414 469152
rect 68278 469140 68284 469152
rect 68336 469140 68342 469192
rect 192018 469140 192024 469192
rect 192076 469180 192082 469192
rect 213086 469180 213092 469192
rect 192076 469152 213092 469180
rect 192076 469140 192082 469152
rect 213086 469140 213092 469152
rect 213144 469140 213150 469192
rect 266354 469140 266360 469192
rect 266412 469180 266418 469192
rect 359734 469180 359740 469192
rect 266412 469152 359740 469180
rect 266412 469140 266418 469152
rect 359734 469140 359740 469152
rect 359792 469140 359798 469192
rect 49602 469072 49608 469124
rect 49660 469112 49666 469124
rect 70578 469112 70584 469124
rect 49660 469084 70584 469112
rect 49660 469072 49666 469084
rect 70578 469072 70584 469084
rect 70636 469072 70642 469124
rect 193398 469072 193404 469124
rect 193456 469112 193462 469124
rect 217594 469112 217600 469124
rect 193456 469084 217600 469112
rect 193456 469072 193462 469084
rect 217594 469072 217600 469084
rect 217652 469072 217658 469124
rect 271966 469072 271972 469124
rect 272024 469112 272030 469124
rect 366174 469112 366180 469124
rect 272024 469084 366180 469112
rect 272024 469072 272030 469084
rect 366174 469072 366180 469084
rect 366232 469072 366238 469124
rect 54938 469004 54944 469056
rect 54996 469044 55002 469056
rect 85666 469044 85672 469056
rect 54996 469016 85672 469044
rect 54996 469004 55002 469016
rect 85666 469004 85672 469016
rect 85724 469004 85730 469056
rect 175274 469004 175280 469056
rect 175332 469044 175338 469056
rect 206646 469044 206652 469056
rect 175332 469016 206652 469044
rect 175332 469004 175338 469016
rect 206646 469004 206652 469016
rect 206704 469004 206710 469056
rect 266538 469004 266544 469056
rect 266596 469044 266602 469056
rect 361206 469044 361212 469056
rect 266596 469016 361212 469044
rect 266596 469004 266602 469016
rect 361206 469004 361212 469016
rect 361264 469004 361270 469056
rect 56042 468936 56048 468988
rect 56100 468976 56106 468988
rect 87138 468976 87144 468988
rect 56100 468948 87144 468976
rect 56100 468936 56106 468948
rect 87138 468936 87144 468948
rect 87196 468936 87202 468988
rect 180886 468936 180892 468988
rect 180944 468976 180950 468988
rect 212350 468976 212356 468988
rect 180944 468948 212356 468976
rect 180944 468936 180950 468948
rect 212350 468936 212356 468948
rect 212408 468936 212414 468988
rect 265158 468936 265164 468988
rect 265216 468976 265222 468988
rect 361114 468976 361120 468988
rect 265216 468948 361120 468976
rect 265216 468936 265222 468948
rect 361114 468936 361120 468948
rect 361172 468936 361178 468988
rect 55030 468868 55036 468920
rect 55088 468908 55094 468920
rect 86954 468908 86960 468920
rect 55088 468880 86960 468908
rect 55088 468868 55094 468880
rect 86954 468868 86960 468880
rect 87012 468868 87018 468920
rect 179414 468868 179420 468920
rect 179472 468908 179478 468920
rect 214742 468908 214748 468920
rect 179472 468880 214748 468908
rect 179472 468868 179478 468880
rect 214742 468868 214748 468880
rect 214800 468868 214806 468920
rect 276014 468868 276020 468920
rect 276072 468908 276078 468920
rect 374362 468908 374368 468920
rect 276072 468880 374368 468908
rect 276072 468868 276078 468880
rect 374362 468868 374368 468880
rect 374420 468868 374426 468920
rect 54846 468800 54852 468852
rect 54904 468840 54910 468852
rect 88518 468840 88524 468852
rect 54904 468812 88524 468840
rect 54904 468800 54910 468812
rect 88518 468800 88524 468812
rect 88576 468800 88582 468852
rect 167178 468800 167184 468852
rect 167236 468840 167242 468852
rect 209130 468840 209136 468852
rect 167236 468812 209136 468840
rect 167236 468800 167242 468812
rect 209130 468800 209136 468812
rect 209188 468800 209194 468852
rect 267734 468800 267740 468852
rect 267792 468840 267798 468852
rect 369026 468840 369032 468852
rect 267792 468812 369032 468840
rect 267792 468800 267798 468812
rect 369026 468800 369032 468812
rect 369084 468800 369090 468852
rect 52086 468732 52092 468784
rect 52144 468772 52150 468784
rect 85574 468772 85580 468784
rect 52144 468744 85580 468772
rect 52144 468732 52150 468744
rect 85574 468732 85580 468744
rect 85632 468732 85638 468784
rect 142338 468732 142344 468784
rect 142396 468772 142402 468784
rect 199010 468772 199016 468784
rect 142396 468744 199016 468772
rect 142396 468732 142402 468744
rect 199010 468732 199016 468744
rect 199068 468732 199074 468784
rect 255314 468732 255320 468784
rect 255372 468772 255378 468784
rect 356790 468772 356796 468784
rect 255372 468744 356796 468772
rect 255372 468732 255378 468744
rect 356790 468732 356796 468744
rect 356848 468732 356854 468784
rect 53466 468664 53472 468716
rect 53524 468704 53530 468716
rect 87046 468704 87052 468716
rect 53524 468676 87052 468704
rect 53524 468664 53530 468676
rect 87046 468664 87052 468676
rect 87104 468664 87110 468716
rect 139394 468664 139400 468716
rect 139452 468704 139458 468716
rect 197262 468704 197268 468716
rect 139452 468676 197268 468704
rect 139452 468664 139458 468676
rect 197262 468664 197268 468676
rect 197320 468664 197326 468716
rect 254026 468664 254032 468716
rect 254084 468704 254090 468716
rect 358538 468704 358544 468716
rect 254084 468676 358544 468704
rect 254084 468664 254090 468676
rect 358538 468664 358544 468676
rect 358596 468664 358602 468716
rect 49326 468596 49332 468648
rect 49384 468636 49390 468648
rect 92566 468636 92572 468648
rect 49384 468608 92572 468636
rect 49384 468596 49390 468608
rect 92566 468596 92572 468608
rect 92624 468596 92630 468648
rect 109034 468596 109040 468648
rect 109092 468636 109098 468648
rect 197722 468636 197728 468648
rect 109092 468608 197728 468636
rect 109092 468596 109098 468608
rect 197722 468596 197728 468608
rect 197780 468596 197786 468648
rect 266446 468596 266452 468648
rect 266504 468636 266510 468648
rect 375282 468636 375288 468648
rect 266504 468608 375288 468636
rect 266504 468596 266510 468608
rect 375282 468596 375288 468608
rect 375340 468596 375346 468648
rect 49234 468528 49240 468580
rect 49292 468568 49298 468580
rect 93946 468568 93952 468580
rect 49292 468540 93952 468568
rect 49292 468528 49298 468540
rect 93946 468528 93952 468540
rect 94004 468528 94010 468580
rect 107746 468528 107752 468580
rect 107804 468568 107810 468580
rect 197630 468568 197636 468580
rect 107804 468540 197636 468568
rect 107804 468528 107810 468540
rect 197630 468528 197636 468540
rect 197688 468528 197694 468580
rect 249978 468528 249984 468580
rect 250036 468568 250042 468580
rect 365162 468568 365168 468580
rect 250036 468540 365168 468568
rect 250036 468528 250042 468540
rect 365162 468528 365168 468540
rect 365220 468528 365226 468580
rect 43346 468460 43352 468512
rect 43404 468500 43410 468512
rect 103514 468500 103520 468512
rect 43404 468472 103520 468500
rect 43404 468460 43410 468472
rect 103514 468460 103520 468472
rect 103572 468460 103578 468512
rect 107654 468460 107660 468512
rect 107712 468500 107718 468512
rect 201678 468500 201684 468512
rect 107712 468472 201684 468500
rect 107712 468460 107718 468472
rect 201678 468460 201684 468472
rect 201736 468460 201742 468512
rect 249886 468460 249892 468512
rect 249944 468500 249950 468512
rect 373350 468500 373356 468512
rect 249944 468472 373356 468500
rect 249944 468460 249950 468472
rect 373350 468460 373356 468472
rect 373408 468460 373414 468512
rect 47670 468392 47676 468444
rect 47728 468432 47734 468444
rect 63586 468432 63592 468444
rect 47728 468404 63592 468432
rect 47728 468392 47734 468404
rect 63586 468392 63592 468404
rect 63644 468392 63650 468444
rect 191926 468392 191932 468444
rect 191984 468432 191990 468444
rect 211614 468432 211620 468444
rect 191984 468404 211620 468432
rect 191984 468392 191990 468404
rect 211614 468392 211620 468404
rect 211672 468392 211678 468444
rect 294046 468392 294052 468444
rect 294104 468432 294110 468444
rect 375742 468432 375748 468444
rect 294104 468404 375748 468432
rect 294104 468392 294110 468404
rect 375742 468392 375748 468404
rect 375800 468392 375806 468444
rect 192110 468324 192116 468376
rect 192168 468364 192174 468376
rect 210050 468364 210056 468376
rect 192168 468336 210056 468364
rect 192168 468324 192174 468336
rect 210050 468324 210056 468336
rect 210108 468324 210114 468376
rect 186314 468256 186320 468308
rect 186372 468296 186378 468308
rect 200850 468296 200856 468308
rect 186372 468268 200856 468296
rect 186372 468256 186378 468268
rect 200850 468256 200856 468268
rect 200908 468256 200914 468308
rect 80698 467780 80704 467832
rect 80756 467820 80762 467832
rect 178034 467820 178040 467832
rect 80756 467792 178040 467820
rect 80756 467780 80762 467792
rect 178034 467780 178040 467792
rect 178092 467780 178098 467832
rect 292666 467576 292672 467628
rect 292724 467616 292730 467628
rect 357986 467616 357992 467628
rect 292724 467588 357992 467616
rect 292724 467576 292730 467588
rect 357986 467576 357992 467588
rect 358044 467576 358050 467628
rect 277486 467508 277492 467560
rect 277544 467548 277550 467560
rect 367646 467548 367652 467560
rect 277544 467520 367652 467548
rect 277544 467508 277550 467520
rect 367646 467508 367652 467520
rect 367704 467508 367710 467560
rect 189166 467440 189172 467492
rect 189224 467480 189230 467492
rect 200758 467480 200764 467492
rect 189224 467452 200764 467480
rect 189224 467440 189230 467452
rect 200758 467440 200764 467452
rect 200816 467440 200822 467492
rect 273254 467440 273260 467492
rect 273312 467480 273318 467492
rect 363506 467480 363512 467492
rect 273312 467452 363512 467480
rect 273312 467440 273318 467452
rect 363506 467440 363512 467452
rect 363564 467440 363570 467492
rect 189074 467372 189080 467424
rect 189132 467412 189138 467424
rect 202506 467412 202512 467424
rect 189132 467384 202512 467412
rect 189132 467372 189138 467384
rect 202506 467372 202512 467384
rect 202564 467372 202570 467424
rect 256694 467372 256700 467424
rect 256752 467412 256758 467424
rect 361022 467412 361028 467424
rect 256752 467384 361028 467412
rect 256752 467372 256758 467384
rect 361022 467372 361028 467384
rect 361080 467372 361086 467424
rect 44082 467304 44088 467356
rect 44140 467344 44146 467356
rect 70486 467344 70492 467356
rect 44140 467316 70492 467344
rect 44140 467304 44146 467316
rect 70486 467304 70492 467316
rect 70544 467304 70550 467356
rect 184934 467304 184940 467356
rect 184992 467344 184998 467356
rect 212166 467344 212172 467356
rect 184992 467316 212172 467344
rect 184992 467304 184998 467316
rect 212166 467304 212172 467316
rect 212224 467304 212230 467356
rect 251266 467304 251272 467356
rect 251324 467344 251330 467356
rect 365254 467344 365260 467356
rect 251324 467316 365260 467344
rect 251324 467304 251330 467316
rect 365254 467304 365260 467316
rect 365312 467304 365318 467356
rect 42242 467236 42248 467288
rect 42300 467276 42306 467288
rect 73798 467276 73804 467288
rect 42300 467248 73804 467276
rect 42300 467236 42306 467248
rect 73798 467236 73804 467248
rect 73856 467236 73862 467288
rect 180150 467236 180156 467288
rect 180208 467276 180214 467288
rect 218054 467276 218060 467288
rect 180208 467248 218060 467276
rect 180208 467236 180214 467248
rect 218054 467236 218060 467248
rect 218112 467236 218118 467288
rect 260834 467236 260840 467288
rect 260892 467276 260898 467288
rect 376294 467276 376300 467288
rect 260892 467248 376300 467276
rect 260892 467236 260898 467248
rect 376294 467236 376300 467248
rect 376352 467236 376358 467288
rect 41322 467168 41328 467220
rect 41380 467208 41386 467220
rect 93854 467208 93860 467220
rect 41380 467180 93860 467208
rect 41380 467168 41386 467180
rect 93854 467168 93860 467180
rect 93912 467168 93918 467220
rect 164234 467168 164240 467220
rect 164292 467208 164298 467220
rect 218882 467208 218888 467220
rect 164292 467180 218888 467208
rect 164292 467168 164298 467180
rect 218882 467168 218888 467180
rect 218940 467168 218946 467220
rect 258074 467168 258080 467220
rect 258132 467208 258138 467220
rect 373626 467208 373632 467220
rect 258132 467180 373632 467208
rect 258132 467168 258138 467180
rect 373626 467168 373632 467180
rect 373684 467168 373690 467220
rect 47946 467100 47952 467152
rect 48004 467140 48010 467152
rect 106458 467140 106464 467152
rect 48004 467112 106464 467140
rect 48004 467100 48010 467112
rect 106458 467100 106464 467112
rect 106516 467100 106522 467152
rect 151814 467100 151820 467152
rect 151872 467140 151878 467152
rect 210418 467140 210424 467152
rect 151872 467112 210424 467140
rect 151872 467100 151878 467112
rect 210418 467100 210424 467112
rect 210476 467100 210482 467152
rect 251174 467100 251180 467152
rect 251232 467140 251238 467152
rect 366910 467140 366916 467152
rect 251232 467112 366916 467140
rect 251232 467100 251238 467112
rect 366910 467100 366916 467112
rect 366968 467100 366974 467152
rect 339402 466556 339408 466608
rect 339460 466596 339466 466608
rect 361574 466596 361580 466608
rect 339460 466568 361580 466596
rect 339460 466556 339466 466568
rect 361574 466556 361580 466568
rect 361632 466596 361638 466608
rect 498470 466596 498476 466608
rect 361632 466568 498476 466596
rect 361632 466556 361638 466568
rect 498470 466556 498476 466568
rect 498528 466596 498534 466608
rect 517882 466596 517888 466608
rect 498528 466568 517888 466596
rect 498528 466556 498534 466568
rect 517882 466556 517888 466568
rect 517940 466556 517946 466608
rect 178034 466488 178040 466540
rect 178092 466528 178098 466540
rect 178092 466500 209774 466528
rect 178092 466488 178098 466500
rect 190914 466420 190920 466472
rect 190972 466460 190978 466472
rect 207014 466460 207020 466472
rect 190972 466432 207020 466460
rect 190972 466420 190978 466432
rect 207014 466420 207020 466432
rect 207072 466420 207078 466472
rect 209746 466460 209774 466500
rect 218054 466488 218060 466540
rect 218112 466528 218118 466540
rect 218238 466528 218244 466540
rect 218112 466500 218244 466528
rect 218112 466488 218118 466500
rect 218238 466488 218244 466500
rect 218296 466528 218302 466540
rect 339770 466528 339776 466540
rect 218296 466500 339776 466528
rect 218296 466488 218302 466500
rect 339770 466488 339776 466500
rect 339828 466528 339834 466540
rect 356974 466528 356980 466540
rect 339828 466500 356980 466528
rect 339828 466488 339834 466500
rect 356974 466488 356980 466500
rect 357032 466528 357038 466540
rect 499758 466528 499764 466540
rect 357032 466500 499764 466528
rect 357032 466488 357038 466500
rect 499758 466488 499764 466500
rect 499816 466528 499822 466540
rect 499816 466500 509234 466528
rect 499816 466488 499822 466500
rect 212810 466460 212816 466472
rect 209746 466432 212816 466460
rect 212810 466420 212816 466432
rect 212868 466460 212874 466472
rect 338482 466460 338488 466472
rect 212868 466432 338488 466460
rect 212868 466420 212874 466432
rect 338482 466420 338488 466432
rect 338540 466460 338546 466472
rect 339402 466460 339408 466472
rect 338540 466432 339408 466460
rect 338540 466420 338546 466432
rect 339402 466420 339408 466432
rect 339460 466420 339466 466472
rect 350994 466420 351000 466472
rect 351052 466460 351058 466472
rect 362954 466460 362960 466472
rect 351052 466432 362960 466460
rect 351052 466420 351058 466432
rect 362954 466420 362960 466432
rect 363012 466420 363018 466472
rect 509206 466460 509234 466500
rect 510890 466488 510896 466540
rect 510948 466528 510954 466540
rect 517514 466528 517520 466540
rect 510948 466500 517520 466528
rect 510948 466488 510954 466500
rect 517514 466488 517520 466500
rect 517572 466488 517578 466540
rect 517790 466460 517796 466472
rect 509206 466432 517796 466460
rect 517790 466420 517796 466432
rect 517848 466420 517854 466472
rect 51994 466352 52000 466404
rect 52052 466392 52058 466404
rect 75914 466392 75920 466404
rect 52052 466364 75920 466392
rect 52052 466352 52058 466364
rect 75914 466352 75920 466364
rect 75972 466352 75978 466404
rect 182174 466352 182180 466404
rect 182232 466392 182238 466404
rect 202414 466392 202420 466404
rect 182232 466364 202420 466392
rect 182232 466352 182238 466364
rect 202414 466352 202420 466364
rect 202472 466352 202478 466404
rect 213822 466352 213828 466404
rect 213880 466392 213886 466404
rect 220998 466392 221004 466404
rect 213880 466364 221004 466392
rect 213880 466352 213886 466364
rect 220998 466352 221004 466364
rect 221056 466352 221062 466404
rect 264974 466352 264980 466404
rect 265032 466392 265038 466404
rect 368198 466392 368204 466404
rect 265032 466364 368204 466392
rect 265032 466352 265038 466364
rect 368198 466352 368204 466364
rect 368256 466352 368262 466404
rect 55674 466284 55680 466336
rect 55732 466324 55738 466336
rect 77478 466324 77484 466336
rect 55732 466296 77484 466324
rect 55732 466284 55738 466296
rect 77478 466284 77484 466296
rect 77536 466284 77542 466336
rect 187694 466284 187700 466336
rect 187752 466324 187758 466336
rect 211522 466324 211528 466336
rect 187752 466296 211528 466324
rect 187752 466284 187758 466296
rect 211522 466284 211528 466296
rect 211580 466284 211586 466336
rect 269114 466284 269120 466336
rect 269172 466324 269178 466336
rect 372522 466324 372528 466336
rect 269172 466296 372528 466324
rect 269172 466284 269178 466296
rect 372522 466284 372528 466296
rect 372580 466284 372586 466336
rect 191834 466216 191840 466268
rect 191892 466256 191898 466268
rect 215846 466256 215852 466268
rect 191892 466228 215852 466256
rect 191892 466216 191898 466228
rect 215846 466216 215852 466228
rect 215904 466216 215910 466268
rect 262214 466216 262220 466268
rect 262272 466256 262278 466268
rect 379054 466256 379060 466268
rect 262272 466228 379060 466256
rect 262272 466216 262278 466228
rect 379054 466216 379060 466228
rect 379112 466216 379118 466268
rect 54386 466148 54392 466200
rect 54444 466188 54450 466200
rect 62114 466188 62120 466200
rect 54444 466160 62120 466188
rect 54444 466148 54450 466160
rect 62114 466148 62120 466160
rect 62172 466148 62178 466200
rect 180794 466148 180800 466200
rect 180852 466188 180858 466200
rect 206738 466188 206744 466200
rect 180852 466160 206744 466188
rect 180852 466148 180858 466160
rect 206738 466148 206744 466160
rect 206796 466148 206802 466200
rect 249794 466148 249800 466200
rect 249852 466188 249858 466200
rect 367922 466188 367928 466200
rect 249852 466160 367928 466188
rect 249852 466148 249858 466160
rect 367922 466148 367928 466160
rect 367980 466148 367986 466200
rect 59262 466080 59268 466132
rect 59320 466120 59326 466132
rect 67634 466120 67640 466132
rect 59320 466092 67640 466120
rect 59320 466080 59326 466092
rect 67634 466080 67640 466092
rect 67692 466080 67698 466132
rect 173986 466080 173992 466132
rect 174044 466120 174050 466132
rect 203794 466120 203800 466132
rect 174044 466092 203800 466120
rect 174044 466080 174050 466092
rect 203794 466080 203800 466092
rect 203852 466080 203858 466132
rect 248506 466080 248512 466132
rect 248564 466120 248570 466132
rect 370682 466120 370688 466132
rect 248564 466092 370688 466120
rect 248564 466080 248570 466092
rect 370682 466080 370688 466092
rect 370740 466080 370746 466132
rect 54294 466012 54300 466064
rect 54352 466052 54358 466064
rect 63494 466052 63500 466064
rect 54352 466024 63500 466052
rect 54352 466012 54358 466024
rect 63494 466012 63500 466024
rect 63552 466012 63558 466064
rect 176654 466012 176660 466064
rect 176712 466052 176718 466064
rect 209406 466052 209412 466064
rect 176712 466024 209412 466052
rect 176712 466012 176718 466024
rect 209406 466012 209412 466024
rect 209464 466012 209470 466064
rect 248414 466012 248420 466064
rect 248472 466052 248478 466064
rect 372154 466052 372160 466064
rect 248472 466024 372160 466052
rect 248472 466012 248478 466024
rect 372154 466012 372160 466024
rect 372212 466012 372218 466064
rect 43254 465944 43260 465996
rect 43312 465984 43318 465996
rect 60826 465984 60832 465996
rect 43312 465956 60832 465984
rect 43312 465944 43318 465956
rect 60826 465944 60832 465956
rect 60884 465944 60890 465996
rect 164878 465944 164884 465996
rect 164936 465984 164942 465996
rect 200298 465984 200304 465996
rect 164936 465956 200304 465984
rect 164936 465944 164942 465956
rect 200298 465944 200304 465956
rect 200356 465944 200362 465996
rect 253934 465944 253940 465996
rect 253992 465984 253998 465996
rect 379146 465984 379152 465996
rect 253992 465956 379152 465984
rect 253992 465944 253998 465956
rect 379146 465944 379152 465956
rect 379204 465944 379210 465996
rect 52270 465876 52276 465928
rect 52328 465916 52334 465928
rect 70394 465916 70400 465928
rect 52328 465888 70400 465916
rect 52328 465876 52334 465888
rect 70394 465876 70400 465888
rect 70452 465876 70458 465928
rect 173894 465876 173900 465928
rect 173952 465916 173958 465928
rect 214834 465916 214840 465928
rect 173952 465888 214840 465916
rect 173952 465876 173958 465888
rect 214834 465876 214840 465888
rect 214892 465876 214898 465928
rect 241514 465876 241520 465928
rect 241572 465916 241578 465928
rect 367830 465916 367836 465928
rect 241572 465888 367836 465916
rect 241572 465876 241578 465888
rect 367830 465876 367836 465888
rect 367888 465876 367894 465928
rect 42150 465808 42156 465860
rect 42208 465848 42214 465860
rect 60734 465848 60740 465860
rect 42208 465820 60740 465848
rect 42208 465808 42214 465820
rect 60734 465808 60740 465820
rect 60792 465808 60798 465860
rect 140774 465808 140780 465860
rect 140832 465848 140838 465860
rect 203242 465848 203248 465860
rect 140832 465820 203248 465848
rect 140832 465808 140838 465820
rect 203242 465808 203248 465820
rect 203300 465808 203306 465860
rect 244274 465808 244280 465860
rect 244332 465848 244338 465860
rect 370590 465848 370596 465860
rect 244332 465820 370596 465848
rect 244332 465808 244338 465820
rect 370590 465808 370596 465820
rect 370648 465808 370654 465860
rect 51442 465740 51448 465792
rect 51500 465780 51506 465792
rect 52178 465780 52184 465792
rect 51500 465752 52184 465780
rect 51500 465740 51506 465752
rect 52178 465740 52184 465752
rect 52236 465740 52242 465792
rect 53742 465740 53748 465792
rect 53800 465780 53806 465792
rect 74718 465780 74724 465792
rect 53800 465752 74724 465780
rect 53800 465740 53806 465752
rect 74718 465740 74724 465752
rect 74776 465740 74782 465792
rect 142246 465740 142252 465792
rect 142304 465780 142310 465792
rect 207382 465780 207388 465792
rect 142304 465752 207388 465780
rect 142304 465740 142310 465752
rect 207382 465740 207388 465752
rect 207440 465740 207446 465792
rect 235994 465740 236000 465792
rect 236052 465780 236058 465792
rect 363782 465780 363788 465792
rect 236052 465752 363788 465780
rect 236052 465740 236058 465752
rect 363782 465740 363788 465752
rect 363840 465740 363846 465792
rect 42702 465672 42708 465724
rect 42760 465712 42766 465724
rect 66346 465712 66352 465724
rect 42760 465684 66352 465712
rect 42760 465672 42766 465684
rect 66346 465672 66352 465684
rect 66404 465672 66410 465724
rect 72418 465672 72424 465724
rect 72476 465712 72482 465724
rect 198918 465712 198924 465724
rect 72476 465684 198924 465712
rect 72476 465672 72482 465684
rect 198918 465672 198924 465684
rect 198976 465672 198982 465724
rect 209682 465672 209688 465724
rect 209740 465712 209746 465724
rect 220906 465712 220912 465724
rect 209740 465684 220912 465712
rect 209740 465672 209746 465684
rect 220906 465672 220912 465684
rect 220964 465672 220970 465724
rect 242894 465672 242900 465724
rect 242952 465712 242958 465724
rect 374730 465712 374736 465724
rect 242952 465684 374736 465712
rect 242952 465672 242958 465684
rect 374730 465672 374736 465684
rect 374788 465672 374794 465724
rect 190546 465604 190552 465656
rect 190604 465644 190610 465656
rect 199470 465644 199476 465656
rect 190604 465616 199476 465644
rect 190604 465604 190610 465616
rect 199470 465604 199476 465616
rect 199528 465604 199534 465656
rect 212994 465644 213000 465656
rect 199580 465616 213000 465644
rect 194594 465536 194600 465588
rect 194652 465576 194658 465588
rect 199580 465576 199608 465616
rect 212994 465604 213000 465616
rect 213052 465604 213058 465656
rect 277394 465604 277400 465656
rect 277452 465644 277458 465656
rect 364702 465644 364708 465656
rect 277452 465616 364708 465644
rect 277452 465604 277458 465616
rect 364702 465604 364708 465616
rect 364760 465604 364766 465656
rect 194652 465548 199608 465576
rect 194652 465536 194658 465548
rect 285674 465536 285680 465588
rect 285732 465576 285738 465588
rect 357894 465576 357900 465588
rect 285732 465548 357900 465576
rect 285732 465536 285738 465548
rect 357894 465536 357900 465548
rect 357952 465536 357958 465588
rect 193306 465468 193312 465520
rect 193364 465508 193370 465520
rect 203886 465508 203892 465520
rect 193364 465480 203892 465508
rect 193364 465468 193370 465480
rect 203886 465468 203892 465480
rect 203944 465468 203950 465520
rect 198918 465060 198924 465112
rect 198976 465100 198982 465112
rect 358814 465100 358820 465112
rect 198976 465072 358820 465100
rect 198976 465060 198982 465072
rect 358814 465060 358820 465072
rect 358872 465100 358878 465112
rect 518894 465100 518900 465112
rect 358872 465072 518900 465100
rect 358872 465060 358878 465072
rect 518894 465060 518900 465072
rect 518952 465060 518958 465112
rect 51350 464992 51356 465044
rect 51408 465032 51414 465044
rect 51994 465032 52000 465044
rect 51408 465004 52000 465032
rect 51408 464992 51414 465004
rect 51994 464992 52000 465004
rect 52052 464992 52058 465044
rect 197170 464992 197176 465044
rect 197228 465032 197234 465044
rect 200574 465032 200580 465044
rect 197228 465004 200580 465032
rect 197228 464992 197234 465004
rect 200574 464992 200580 465004
rect 200632 464992 200638 465044
rect 207474 464992 207480 465044
rect 207532 465032 207538 465044
rect 207934 465032 207940 465044
rect 207532 465004 207940 465032
rect 207532 464992 207538 465004
rect 207934 464992 207940 465004
rect 207992 464992 207998 465044
rect 190454 464720 190460 464772
rect 190512 464760 190518 464772
rect 208762 464760 208768 464772
rect 190512 464732 208768 464760
rect 190512 464720 190518 464732
rect 208762 464720 208768 464732
rect 208820 464720 208826 464772
rect 59078 464652 59084 464704
rect 59136 464692 59142 464704
rect 89898 464692 89904 464704
rect 59136 464664 89904 464692
rect 59136 464652 59142 464664
rect 89898 464652 89904 464664
rect 89956 464652 89962 464704
rect 183646 464652 183652 464704
rect 183704 464692 183710 464704
rect 205266 464692 205272 464704
rect 183704 464664 205272 464692
rect 183704 464652 183710 464664
rect 205266 464652 205272 464664
rect 205324 464652 205330 464704
rect 58986 464584 58992 464636
rect 59044 464624 59050 464636
rect 92474 464624 92480 464636
rect 59044 464596 92480 464624
rect 59044 464584 59050 464596
rect 92474 464584 92480 464596
rect 92532 464584 92538 464636
rect 183554 464584 183560 464636
rect 183612 464624 183618 464636
rect 207842 464624 207848 464636
rect 183612 464596 207848 464624
rect 183612 464584 183618 464596
rect 207842 464584 207848 464596
rect 207900 464584 207906 464636
rect 55858 464516 55864 464568
rect 55916 464556 55922 464568
rect 102318 464556 102324 464568
rect 55916 464528 102324 464556
rect 55916 464516 55922 464528
rect 102318 464516 102324 464528
rect 102376 464516 102382 464568
rect 193214 464516 193220 464568
rect 193272 464556 193278 464568
rect 217778 464556 217784 464568
rect 193272 464528 217784 464556
rect 193272 464516 193278 464528
rect 217778 464516 217784 464528
rect 217836 464516 217842 464568
rect 52914 464448 52920 464500
rect 52972 464488 52978 464500
rect 121454 464488 121460 464500
rect 52972 464460 121460 464488
rect 52972 464448 52978 464460
rect 121454 464448 121460 464460
rect 121512 464448 121518 464500
rect 126974 464448 126980 464500
rect 127032 464488 127038 464500
rect 197814 464488 197820 464500
rect 127032 464460 197820 464488
rect 127032 464448 127038 464460
rect 197814 464448 197820 464460
rect 197872 464448 197878 464500
rect 57054 464380 57060 464432
rect 57112 464420 57118 464432
rect 128354 464420 128360 464432
rect 57112 464392 128360 464420
rect 57112 464380 57118 464392
rect 128354 464380 128360 464392
rect 128412 464380 128418 464432
rect 142154 464380 142160 464432
rect 142212 464420 142218 464432
rect 197998 464420 198004 464432
rect 142212 464392 198004 464420
rect 142212 464380 142218 464392
rect 197998 464380 198004 464392
rect 198056 464380 198062 464432
rect 293954 464380 293960 464432
rect 294012 464420 294018 464432
rect 375006 464420 375012 464432
rect 294012 464392 375012 464420
rect 294012 464380 294018 464392
rect 375006 464380 375012 464392
rect 375064 464380 375070 464432
rect 55950 464312 55956 464364
rect 56008 464352 56014 464364
rect 130010 464352 130016 464364
rect 56008 464324 130016 464352
rect 56008 464312 56014 464324
rect 130010 464312 130016 464324
rect 130068 464312 130074 464364
rect 136634 464312 136640 464364
rect 136692 464352 136698 464364
rect 199286 464352 199292 464364
rect 136692 464324 199292 464352
rect 136692 464312 136698 464324
rect 199286 464312 199292 464324
rect 199344 464312 199350 464364
rect 271874 464312 271880 464364
rect 271932 464352 271938 464364
rect 371786 464352 371792 464364
rect 271932 464324 371792 464352
rect 271932 464312 271938 464324
rect 371786 464312 371792 464324
rect 371844 464312 371850 464364
rect 46014 464244 46020 464296
rect 46072 464284 46078 464296
rect 207934 464284 207940 464296
rect 46072 464256 207940 464284
rect 46072 464244 46078 464256
rect 207934 464244 207940 464256
rect 207992 464244 207998 464296
rect 207934 422900 207940 422952
rect 207992 422940 207998 422952
rect 217962 422940 217968 422952
rect 207992 422912 217968 422940
rect 207992 422900 207998 422912
rect 217962 422900 217968 422912
rect 218020 422900 218026 422952
rect 55674 418208 55680 418260
rect 55732 418248 55738 418260
rect 57146 418248 57152 418260
rect 55732 418220 57152 418248
rect 55732 418208 55738 418220
rect 57146 418208 57152 418220
rect 57204 418208 57210 418260
rect 55766 418140 55772 418192
rect 55824 418180 55830 418192
rect 56870 418180 56876 418192
rect 55824 418152 56876 418180
rect 55824 418140 55830 418152
rect 56870 418140 56876 418152
rect 56928 418140 56934 418192
rect 46014 418072 46020 418124
rect 46072 418112 46078 418124
rect 56962 418112 56968 418124
rect 46072 418084 56968 418112
rect 46072 418072 46078 418084
rect 56962 418072 56968 418084
rect 57020 418072 57026 418124
rect 207198 417460 207204 417512
rect 207256 417500 207262 417512
rect 216674 417500 216680 417512
rect 207256 417472 216680 417500
rect 207256 417460 207262 417472
rect 216674 417460 216680 417472
rect 216732 417460 216738 417512
rect 206830 417392 206836 417444
rect 206888 417432 206894 417444
rect 219618 417432 219624 417444
rect 206888 417404 219624 417432
rect 206888 417392 206894 417404
rect 219618 417392 219624 417404
rect 219676 417392 219682 417444
rect 357894 417392 357900 417444
rect 357952 417432 357958 417444
rect 376938 417432 376944 417444
rect 357952 417404 376944 417432
rect 357952 417392 357958 417404
rect 376938 417392 376944 417404
rect 376996 417392 377002 417444
rect 44634 416780 44640 416832
rect 44692 416820 44698 416832
rect 57882 416820 57888 416832
rect 44692 416792 57888 416820
rect 44692 416780 44698 416792
rect 57882 416780 57888 416792
rect 57940 416780 57946 416832
rect 205818 416712 205824 416764
rect 205876 416752 205882 416764
rect 207934 416752 207940 416764
rect 205876 416724 207940 416752
rect 205876 416712 205882 416724
rect 207934 416712 207940 416724
rect 207992 416712 207998 416764
rect 55674 415352 55680 415404
rect 55732 415392 55738 415404
rect 57054 415392 57060 415404
rect 55732 415364 57060 415392
rect 55732 415352 55738 415364
rect 57054 415352 57060 415364
rect 57112 415352 57118 415404
rect 57146 415352 57152 415404
rect 57204 415392 57210 415404
rect 58434 415392 58440 415404
rect 57204 415364 58440 415392
rect 57204 415352 57210 415364
rect 58434 415352 58440 415364
rect 58492 415352 58498 415404
rect 207934 414808 207940 414860
rect 207992 414848 207998 414860
rect 217134 414848 217140 414860
rect 207992 414820 217140 414848
rect 207992 414808 207998 414820
rect 217134 414808 217140 414820
rect 217192 414808 217198 414860
rect 208118 414740 208124 414792
rect 208176 414780 208182 414792
rect 216858 414780 216864 414792
rect 208176 414752 216864 414780
rect 208176 414740 208182 414752
rect 216858 414740 216864 414752
rect 216916 414740 216922 414792
rect 206922 414672 206928 414724
rect 206980 414712 206986 414724
rect 216766 414712 216772 414724
rect 206980 414684 216772 414712
rect 206980 414672 206986 414684
rect 216766 414672 216772 414684
rect 216824 414672 216830 414724
rect 359826 414672 359832 414724
rect 359884 414712 359890 414724
rect 377674 414712 377680 414724
rect 359884 414684 377680 414712
rect 359884 414672 359890 414684
rect 377674 414672 377680 414684
rect 377732 414672 377738 414724
rect 47578 413992 47584 414044
rect 47636 414032 47642 414044
rect 57882 414032 57888 414044
rect 47636 414004 57888 414032
rect 47636 413992 47642 414004
rect 57882 413992 57888 414004
rect 57940 413992 57946 414044
rect 57238 413924 57244 413976
rect 57296 413964 57302 413976
rect 58434 413964 58440 413976
rect 57296 413936 58440 413964
rect 57296 413924 57302 413936
rect 58434 413924 58440 413936
rect 58492 413924 58498 413976
rect 205726 413244 205732 413296
rect 205784 413284 205790 413296
rect 216858 413284 216864 413296
rect 205784 413256 216864 413284
rect 205784 413244 205790 413256
rect 216858 413244 216864 413256
rect 216916 413244 216922 413296
rect 47486 412632 47492 412684
rect 47544 412672 47550 412684
rect 57882 412672 57888 412684
rect 47544 412644 57888 412672
rect 47544 412632 47550 412644
rect 57882 412632 57888 412644
rect 57940 412632 57946 412684
rect 204438 411884 204444 411936
rect 204496 411924 204502 411936
rect 205726 411924 205732 411936
rect 204496 411896 205732 411924
rect 204496 411884 204502 411896
rect 205726 411884 205732 411896
rect 205784 411884 205790 411936
rect 358078 411884 358084 411936
rect 358136 411924 358142 411936
rect 377030 411924 377036 411936
rect 358136 411896 377036 411924
rect 358136 411884 358142 411896
rect 377030 411884 377036 411896
rect 377088 411884 377094 411936
rect 48222 411272 48228 411324
rect 48280 411312 48286 411324
rect 57882 411312 57888 411324
rect 48280 411284 57888 411312
rect 48280 411272 48286 411284
rect 57882 411272 57888 411284
rect 57940 411272 57946 411324
rect 217778 411272 217784 411324
rect 217836 411312 217842 411324
rect 219250 411312 219256 411324
rect 217836 411284 219256 411312
rect 217836 411272 217842 411284
rect 219250 411272 219256 411284
rect 219308 411272 219314 411324
rect 3326 411204 3332 411256
rect 3384 411244 3390 411256
rect 15838 411244 15844 411256
rect 3384 411216 15844 411244
rect 3384 411204 3390 411216
rect 15838 411204 15844 411216
rect 15896 411204 15902 411256
rect 205726 410524 205732 410576
rect 205784 410564 205790 410576
rect 216766 410564 216772 410576
rect 205784 410536 216772 410564
rect 205784 410524 205790 410536
rect 216766 410524 216772 410536
rect 216824 410564 216830 410576
rect 216950 410564 216956 410576
rect 216824 410536 216956 410564
rect 216824 410524 216830 410536
rect 216950 410524 216956 410536
rect 217008 410524 217014 410576
rect 360010 410524 360016 410576
rect 360068 410564 360074 410576
rect 377030 410564 377036 410576
rect 360068 410536 377036 410564
rect 360068 410524 360074 410536
rect 377030 410524 377036 410536
rect 377088 410564 377094 410576
rect 377490 410564 377496 410576
rect 377088 410536 377496 410564
rect 377088 410524 377094 410536
rect 377490 410524 377496 410536
rect 377548 410524 377554 410576
rect 50246 409844 50252 409896
rect 50304 409884 50310 409896
rect 57882 409884 57888 409896
rect 50304 409856 57888 409884
rect 50304 409844 50310 409856
rect 57882 409844 57888 409856
rect 57940 409844 57946 409896
rect 377950 409844 377956 409896
rect 378008 409884 378014 409896
rect 379422 409884 379428 409896
rect 378008 409856 379428 409884
rect 378008 409844 378014 409856
rect 379422 409844 379428 409856
rect 379480 409844 379486 409896
rect 359918 409096 359924 409148
rect 359976 409136 359982 409148
rect 377398 409136 377404 409148
rect 359976 409108 377404 409136
rect 359976 409096 359982 409108
rect 377398 409096 377404 409108
rect 377456 409096 377462 409148
rect 50982 408484 50988 408536
rect 51040 408524 51046 408536
rect 57882 408524 57888 408536
rect 51040 408496 57888 408524
rect 51040 408484 51046 408496
rect 57882 408484 57888 408496
rect 57940 408484 57946 408536
rect 576118 405628 576124 405680
rect 576176 405668 576182 405680
rect 580166 405668 580172 405680
rect 576176 405640 580172 405668
rect 576176 405628 576182 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 199194 398216 199200 398268
rect 199252 398256 199258 398268
rect 199746 398256 199752 398268
rect 199252 398228 199752 398256
rect 199252 398216 199258 398228
rect 199746 398216 199752 398228
rect 199804 398216 199810 398268
rect 198090 397808 198096 397860
rect 198148 397848 198154 397860
rect 199102 397848 199108 397860
rect 198148 397820 199108 397848
rect 198148 397808 198154 397820
rect 199102 397808 199108 397820
rect 199160 397808 199166 397860
rect 520918 396720 520924 396772
rect 520976 396760 520982 396772
rect 580350 396760 580356 396772
rect 520976 396732 580356 396760
rect 520976 396720 520982 396732
rect 580350 396720 580356 396732
rect 580408 396720 580414 396772
rect 44726 391892 44732 391944
rect 44784 391932 44790 391944
rect 57054 391932 57060 391944
rect 44784 391904 57060 391932
rect 44784 391892 44790 391904
rect 57054 391892 57060 391904
rect 57112 391892 57118 391944
rect 209590 391892 209596 391944
rect 209648 391932 209654 391944
rect 216674 391932 216680 391944
rect 209648 391904 216680 391932
rect 209648 391892 209654 391904
rect 216674 391892 216680 391904
rect 216732 391892 216738 391944
rect 359642 391892 359648 391944
rect 359700 391932 359706 391944
rect 376938 391932 376944 391944
rect 359700 391904 376944 391932
rect 359700 391892 359706 391904
rect 376938 391892 376944 391904
rect 376996 391892 377002 391944
rect 207014 390464 207020 390516
rect 207072 390504 207078 390516
rect 216674 390504 216680 390516
rect 207072 390476 216680 390504
rect 207072 390464 207078 390476
rect 216674 390464 216680 390476
rect 216732 390464 216738 390516
rect 358078 390464 358084 390516
rect 358136 390504 358142 390516
rect 362954 390504 362960 390516
rect 358136 390476 362960 390504
rect 358136 390464 358142 390476
rect 362954 390464 362960 390476
rect 363012 390504 363018 390516
rect 376938 390504 376944 390516
rect 363012 390476 376944 390504
rect 363012 390464 363018 390476
rect 376938 390464 376944 390476
rect 376996 390464 377002 390516
rect 57514 389376 57520 389428
rect 57572 389376 57578 389428
rect 57532 389280 57560 389376
rect 57532 389252 57652 389280
rect 52362 389104 52368 389156
rect 52420 389144 52426 389156
rect 57238 389144 57244 389156
rect 52420 389116 57244 389144
rect 52420 389104 52426 389116
rect 57238 389104 57244 389116
rect 57296 389144 57302 389156
rect 57514 389144 57520 389156
rect 57296 389116 57520 389144
rect 57296 389104 57302 389116
rect 57514 389104 57520 389116
rect 57572 389104 57578 389156
rect 46106 389036 46112 389088
rect 46164 389076 46170 389088
rect 57054 389076 57060 389088
rect 46164 389048 57060 389076
rect 46164 389036 46170 389048
rect 57054 389036 57060 389048
rect 57112 389036 57118 389088
rect 57514 388968 57520 389020
rect 57572 389008 57578 389020
rect 57624 389008 57652 389252
rect 206278 389172 206284 389224
rect 206336 389212 206342 389224
rect 207014 389212 207020 389224
rect 206336 389184 207020 389212
rect 206336 389172 206342 389184
rect 207014 389172 207020 389184
rect 207072 389172 207078 389224
rect 200758 389104 200764 389156
rect 200816 389144 200822 389156
rect 216674 389144 216680 389156
rect 200816 389116 216680 389144
rect 200816 389104 200822 389116
rect 216674 389104 216680 389116
rect 216732 389104 216738 389156
rect 359734 389104 359740 389156
rect 359792 389144 359798 389156
rect 376938 389144 376944 389156
rect 359792 389116 376944 389144
rect 359792 389104 359798 389116
rect 376938 389104 376944 389116
rect 376996 389104 377002 389156
rect 57572 388980 57652 389008
rect 57572 388968 57578 388980
rect 57330 387744 57336 387796
rect 57388 387784 57394 387796
rect 58618 387784 58624 387796
rect 57388 387756 58624 387784
rect 57388 387744 57394 387756
rect 58618 387744 58624 387756
rect 58676 387744 58682 387796
rect 58526 387676 58532 387728
rect 58584 387716 58590 387728
rect 59354 387716 59360 387728
rect 58584 387688 59360 387716
rect 58584 387676 58590 387688
rect 59354 387676 59360 387688
rect 59412 387676 59418 387728
rect 57882 387132 57888 387184
rect 57940 387172 57946 387184
rect 59722 387172 59728 387184
rect 57940 387144 59728 387172
rect 57940 387132 57946 387144
rect 59722 387132 59728 387144
rect 59780 387132 59786 387184
rect 56962 386316 56968 386368
rect 57020 386356 57026 386368
rect 59722 386356 59728 386368
rect 57020 386328 59728 386356
rect 57020 386316 57026 386328
rect 59722 386316 59728 386328
rect 59780 386316 59786 386368
rect 369026 385704 369032 385756
rect 369084 385744 369090 385756
rect 372798 385744 372804 385756
rect 369084 385716 372804 385744
rect 369084 385704 369090 385716
rect 372798 385704 372804 385716
rect 372856 385704 372862 385756
rect 219526 382372 219532 382424
rect 219584 382412 219590 382424
rect 219894 382412 219900 382424
rect 219584 382384 219900 382412
rect 219584 382372 219590 382384
rect 219894 382372 219900 382384
rect 219952 382372 219958 382424
rect 217410 382236 217416 382288
rect 217468 382276 217474 382288
rect 219526 382276 219532 382288
rect 217468 382248 219532 382276
rect 217468 382236 217474 382248
rect 219526 382236 219532 382248
rect 219584 382236 219590 382288
rect 57422 381624 57428 381676
rect 57480 381664 57486 381676
rect 59538 381664 59544 381676
rect 57480 381636 59544 381664
rect 57480 381624 57486 381636
rect 59538 381624 59544 381636
rect 59596 381624 59602 381676
rect 197170 381488 197176 381540
rect 197228 381528 197234 381540
rect 218238 381528 218244 381540
rect 197228 381500 218244 381528
rect 197228 381488 197234 381500
rect 218238 381488 218244 381500
rect 218296 381488 218302 381540
rect 55674 381012 55680 381064
rect 55732 381052 55738 381064
rect 59446 381052 59452 381064
rect 55732 381024 59452 381052
rect 55732 381012 55738 381024
rect 59446 381012 59452 381024
rect 59504 381012 59510 381064
rect 196526 381012 196532 381064
rect 196584 381052 196590 381064
rect 212810 381052 212816 381064
rect 196584 381024 212816 381052
rect 196584 381012 196590 381024
rect 212810 381012 212816 381024
rect 212868 381012 212874 381064
rect 196986 380944 196992 380996
rect 197044 380984 197050 380996
rect 198182 380984 198188 380996
rect 197044 380956 198188 380984
rect 197044 380944 197050 380956
rect 198182 380944 198188 380956
rect 198240 380944 198246 380996
rect 199470 380944 199476 380996
rect 199528 380984 199534 380996
rect 256050 380984 256056 380996
rect 199528 380956 256056 380984
rect 199528 380944 199534 380956
rect 256050 380944 256056 380956
rect 256108 380944 256114 380996
rect 55858 380876 55864 380928
rect 55916 380916 55922 380928
rect 60090 380916 60096 380928
rect 55916 380888 60096 380916
rect 55916 380876 55922 380888
rect 60090 380876 60096 380888
rect 60148 380876 60154 380928
rect 143534 380876 143540 380928
rect 143592 380916 143598 380928
rect 205910 380916 205916 380928
rect 143592 380888 205916 380916
rect 143592 380876 143598 380888
rect 205910 380876 205916 380888
rect 205968 380876 205974 380928
rect 375190 380876 375196 380928
rect 375248 380916 375254 380928
rect 422846 380916 422852 380928
rect 375248 380888 422852 380916
rect 375248 380876 375254 380888
rect 422846 380876 422852 380888
rect 422904 380876 422910 380928
rect 47486 380808 47492 380860
rect 47544 380848 47550 380860
rect 216858 380848 216864 380860
rect 47544 380820 216864 380848
rect 47544 380808 47550 380820
rect 216858 380808 216864 380820
rect 216916 380808 216922 380860
rect 48222 380740 48228 380792
rect 48280 380780 48286 380792
rect 217318 380780 217324 380792
rect 48280 380752 217324 380780
rect 48280 380740 48286 380752
rect 217318 380740 217324 380752
rect 217376 380740 217382 380792
rect 52914 380672 52920 380724
rect 52972 380712 52978 380724
rect 55858 380712 55864 380724
rect 52972 380684 55864 380712
rect 52972 380672 52978 380684
rect 55858 380672 55864 380684
rect 55916 380672 55922 380724
rect 216950 380712 216956 380724
rect 64846 380684 216956 380712
rect 50246 380604 50252 380656
rect 50304 380644 50310 380656
rect 64846 380644 64874 380684
rect 216950 380672 216956 380684
rect 217008 380672 217014 380724
rect 367554 380672 367560 380724
rect 367612 380712 367618 380724
rect 377950 380712 377956 380724
rect 367612 380684 377956 380712
rect 367612 380672 367618 380684
rect 377950 380672 377956 380684
rect 378008 380672 378014 380724
rect 50304 380616 64874 380644
rect 50304 380604 50310 380616
rect 160922 380604 160928 380656
rect 160980 380644 160986 380656
rect 207382 380644 207388 380656
rect 160980 380616 207388 380644
rect 160980 380604 160986 380616
rect 207382 380604 207388 380616
rect 207440 380604 207446 380656
rect 365530 380604 365536 380656
rect 365588 380644 365594 380656
rect 376662 380644 376668 380656
rect 365588 380616 376668 380644
rect 365588 380604 365594 380616
rect 376662 380604 376668 380616
rect 376720 380604 376726 380656
rect 377214 380604 377220 380656
rect 377272 380644 377278 380656
rect 430942 380644 430948 380656
rect 377272 380616 430948 380644
rect 377272 380604 377278 380616
rect 430942 380604 430948 380616
rect 431000 380604 431006 380656
rect 146018 380536 146024 380588
rect 146076 380576 146082 380588
rect 207290 380576 207296 380588
rect 146076 380548 207296 380576
rect 146076 380536 146082 380548
rect 207290 380536 207296 380548
rect 207348 380536 207354 380588
rect 360654 380536 360660 380588
rect 360712 380576 360718 380588
rect 369854 380576 369860 380588
rect 360712 380548 369860 380576
rect 360712 380536 360718 380548
rect 369854 380536 369860 380548
rect 369912 380536 369918 380588
rect 371786 380536 371792 380588
rect 371844 380576 371850 380588
rect 433610 380576 433616 380588
rect 371844 380548 433616 380576
rect 371844 380536 371850 380548
rect 433610 380536 433616 380548
rect 433668 380536 433674 380588
rect 59722 380468 59728 380520
rect 59780 380508 59786 380520
rect 118418 380508 118424 380520
rect 59780 380480 118424 380508
rect 59780 380468 59786 380480
rect 118418 380468 118424 380480
rect 118476 380468 118482 380520
rect 133506 380468 133512 380520
rect 133564 380508 133570 380520
rect 203150 380508 203156 380520
rect 133564 380480 203156 380508
rect 133564 380468 133570 380480
rect 203150 380468 203156 380480
rect 203208 380468 203214 380520
rect 204346 380468 204352 380520
rect 204404 380508 204410 380520
rect 213638 380508 213644 380520
rect 204404 380480 213644 380508
rect 204404 380468 204410 380480
rect 213638 380468 213644 380480
rect 213696 380468 213702 380520
rect 358630 380468 358636 380520
rect 358688 380508 358694 380520
rect 421098 380508 421104 380520
rect 358688 380480 421104 380508
rect 358688 380468 358694 380480
rect 421098 380468 421104 380480
rect 421156 380468 421162 380520
rect 57882 380400 57888 380452
rect 57940 380440 57946 380452
rect 116026 380440 116032 380452
rect 57940 380412 116032 380440
rect 57940 380400 57946 380412
rect 116026 380400 116032 380412
rect 116084 380400 116090 380452
rect 135898 380400 135904 380452
rect 135956 380440 135962 380452
rect 200574 380440 200580 380452
rect 135956 380412 200580 380440
rect 135956 380400 135962 380412
rect 200574 380400 200580 380412
rect 200632 380400 200638 380452
rect 202966 380400 202972 380452
rect 203024 380440 203030 380452
rect 274634 380440 274640 380452
rect 203024 380412 274640 380440
rect 203024 380400 203030 380412
rect 274634 380400 274640 380412
rect 274692 380400 274698 380452
rect 369670 380400 369676 380452
rect 369728 380440 369734 380452
rect 436002 380440 436008 380452
rect 369728 380412 436008 380440
rect 369728 380400 369734 380412
rect 436002 380400 436008 380412
rect 436060 380400 436066 380452
rect 48774 380332 48780 380384
rect 48832 380372 48838 380384
rect 110966 380372 110972 380384
rect 48832 380344 110972 380372
rect 48832 380332 48838 380344
rect 110966 380332 110972 380344
rect 111024 380332 111030 380384
rect 131022 380332 131028 380384
rect 131080 380372 131086 380384
rect 204622 380372 204628 380384
rect 131080 380344 204628 380372
rect 131080 380332 131086 380344
rect 204622 380332 204628 380344
rect 204680 380332 204686 380384
rect 262858 380332 262864 380384
rect 262916 380372 262922 380384
rect 269758 380372 269764 380384
rect 262916 380344 269764 380372
rect 262916 380332 262922 380344
rect 269758 380332 269764 380344
rect 269816 380332 269822 380384
rect 366174 380332 366180 380384
rect 366232 380372 366238 380384
rect 438486 380372 438492 380384
rect 366232 380344 438492 380372
rect 366232 380332 366238 380344
rect 438486 380332 438492 380344
rect 438544 380332 438550 380384
rect 58434 380264 58440 380316
rect 58492 380304 58498 380316
rect 123478 380304 123484 380316
rect 58492 380276 123484 380304
rect 58492 380264 58498 380276
rect 123478 380264 123484 380276
rect 123536 380264 123542 380316
rect 163406 380264 163412 380316
rect 163464 380304 163470 380316
rect 197998 380304 198004 380316
rect 163464 380276 198004 380304
rect 163464 380264 163470 380276
rect 197998 380264 198004 380276
rect 198056 380264 198062 380316
rect 200114 380264 200120 380316
rect 200172 380304 200178 380316
rect 293954 380304 293960 380316
rect 200172 380276 293960 380304
rect 200172 380264 200178 380276
rect 293954 380264 293960 380276
rect 294012 380264 294018 380316
rect 363506 380264 363512 380316
rect 363564 380304 363570 380316
rect 440878 380304 440884 380316
rect 363564 380276 440884 380304
rect 363564 380264 363570 380276
rect 440878 380264 440884 380276
rect 440936 380264 440942 380316
rect 58618 380196 58624 380248
rect 58676 380236 58682 380248
rect 125962 380236 125968 380248
rect 58676 380208 125968 380236
rect 58676 380196 58682 380208
rect 125962 380196 125968 380208
rect 126020 380196 126026 380248
rect 128354 380196 128360 380248
rect 128412 380236 128418 380248
rect 199286 380236 199292 380248
rect 128412 380208 199292 380236
rect 128412 380196 128418 380208
rect 199286 380196 199292 380208
rect 199344 380196 199350 380248
rect 200206 380196 200212 380248
rect 200264 380236 200270 380248
rect 301498 380236 301504 380248
rect 200264 380208 301504 380236
rect 200264 380196 200270 380208
rect 301498 380196 301504 380208
rect 301556 380196 301562 380248
rect 360746 380196 360752 380248
rect 360804 380236 360810 380248
rect 443454 380236 443460 380248
rect 360804 380208 443460 380236
rect 360804 380196 360810 380208
rect 443454 380196 443460 380208
rect 443512 380196 443518 380248
rect 45002 380128 45008 380180
rect 45060 380168 45066 380180
rect 113542 380168 113548 380180
rect 45060 380140 113548 380168
rect 45060 380128 45066 380140
rect 113542 380128 113548 380140
rect 113600 380128 113606 380180
rect 120994 380128 121000 380180
rect 121052 380168 121058 380180
rect 197906 380168 197912 380180
rect 121052 380140 197912 380168
rect 121052 380128 121058 380140
rect 197906 380128 197912 380140
rect 197964 380128 197970 380180
rect 201586 380128 201592 380180
rect 201644 380168 201650 380180
rect 309042 380168 309048 380180
rect 201644 380140 309048 380168
rect 201644 380128 201650 380140
rect 309042 380128 309048 380140
rect 309100 380128 309106 380180
rect 362862 380128 362868 380180
rect 362920 380168 362926 380180
rect 445938 380168 445944 380180
rect 362920 380140 445944 380168
rect 362920 380128 362926 380140
rect 445938 380128 445944 380140
rect 445996 380128 446002 380180
rect 155954 380060 155960 380112
rect 156012 380100 156018 380112
rect 203242 380100 203248 380112
rect 156012 380072 203248 380100
rect 156012 380060 156018 380072
rect 203242 380060 203248 380072
rect 203300 380060 203306 380112
rect 158530 379992 158536 380044
rect 158588 380032 158594 380044
rect 201862 380032 201868 380044
rect 158588 380004 201868 380032
rect 158588 379992 158594 380004
rect 201862 379992 201868 380004
rect 201920 379992 201926 380044
rect 214926 379992 214932 380044
rect 214984 380032 214990 380044
rect 218054 380032 218060 380044
rect 214984 380004 218060 380032
rect 214984 379992 214990 380004
rect 218054 379992 218060 380004
rect 218112 379992 218118 380044
rect 165982 379924 165988 379976
rect 166040 379964 166046 379976
rect 199010 379964 199016 379976
rect 166040 379936 199016 379964
rect 166040 379924 166046 379936
rect 199010 379924 199016 379936
rect 199068 379924 199074 379976
rect 213730 379924 213736 379976
rect 213788 379964 213794 379976
rect 235994 379964 236000 379976
rect 213788 379936 236000 379964
rect 213788 379924 213794 379936
rect 235994 379924 236000 379936
rect 236052 379924 236058 379976
rect 240042 379924 240048 379976
rect 240100 379964 240106 379976
rect 259454 379964 259460 379976
rect 240100 379936 259460 379964
rect 240100 379924 240106 379936
rect 259454 379924 259460 379936
rect 259512 379924 259518 379976
rect 207106 379856 207112 379908
rect 207164 379896 207170 379908
rect 216490 379896 216496 379908
rect 207164 379868 216496 379896
rect 207164 379856 207170 379868
rect 216490 379856 216496 379868
rect 216548 379896 216554 379908
rect 243078 379896 243084 379908
rect 216548 379868 243084 379896
rect 216548 379856 216554 379868
rect 243078 379856 243084 379868
rect 243136 379856 243142 379908
rect 213638 379788 213644 379840
rect 213696 379828 213702 379840
rect 237098 379828 237104 379840
rect 213696 379800 237104 379828
rect 213696 379788 213702 379800
rect 237098 379788 237104 379800
rect 237156 379788 237162 379840
rect 237374 379788 237380 379840
rect 237432 379828 237438 379840
rect 265250 379828 265256 379840
rect 237432 379800 265256 379828
rect 237432 379788 237438 379800
rect 265250 379788 265256 379800
rect 265308 379788 265314 379840
rect 377398 379788 377404 379840
rect 377456 379828 377462 379840
rect 377950 379828 377956 379840
rect 377456 379800 377956 379828
rect 377456 379788 377462 379800
rect 377950 379788 377956 379800
rect 378008 379828 378014 379840
rect 408678 379828 408684 379840
rect 378008 379800 408684 379828
rect 378008 379788 378014 379800
rect 408678 379788 408684 379800
rect 408736 379788 408742 379840
rect 212626 379720 212632 379772
rect 212684 379760 212690 379772
rect 213914 379760 213920 379772
rect 212684 379732 213920 379760
rect 212684 379720 212690 379732
rect 213914 379720 213920 379732
rect 213972 379760 213978 379772
rect 220814 379760 220820 379772
rect 213972 379732 220820 379760
rect 213972 379720 213978 379732
rect 220814 379720 220820 379732
rect 220872 379720 220878 379772
rect 254486 379760 254492 379772
rect 220924 379732 254492 379760
rect 212718 379652 212724 379704
rect 212776 379692 212782 379704
rect 219434 379692 219440 379704
rect 212776 379664 219440 379692
rect 212776 379652 212782 379664
rect 219434 379652 219440 379664
rect 219492 379692 219498 379704
rect 220924 379692 220952 379732
rect 254486 379720 254492 379732
rect 254544 379720 254550 379772
rect 369854 379720 369860 379772
rect 369912 379760 369918 379772
rect 370958 379760 370964 379772
rect 369912 379732 370964 379760
rect 369912 379720 369918 379732
rect 370958 379720 370964 379732
rect 371016 379760 371022 379772
rect 413462 379760 413468 379772
rect 371016 379732 413468 379760
rect 371016 379720 371022 379732
rect 413462 379720 413468 379732
rect 413520 379720 413526 379772
rect 219492 379664 220952 379692
rect 219492 379652 219498 379664
rect 220998 379652 221004 379704
rect 221056 379692 221062 379704
rect 255866 379692 255872 379704
rect 221056 379664 255872 379692
rect 221056 379652 221062 379664
rect 255866 379652 255872 379664
rect 255924 379652 255930 379704
rect 376478 379652 376484 379704
rect 376536 379692 376542 379704
rect 376662 379692 376668 379704
rect 376536 379664 376668 379692
rect 376536 379652 376542 379664
rect 376662 379652 376668 379664
rect 376720 379692 376726 379704
rect 419442 379692 419448 379704
rect 376720 379664 419448 379692
rect 376720 379652 376726 379664
rect 419442 379652 419448 379664
rect 419500 379652 419506 379704
rect 208118 379584 208124 379636
rect 208176 379624 208182 379636
rect 209498 379624 209504 379636
rect 208176 379596 209504 379624
rect 208176 379584 208182 379596
rect 209498 379584 209504 379596
rect 209556 379584 209562 379636
rect 216950 379584 216956 379636
rect 217008 379624 217014 379636
rect 217778 379624 217784 379636
rect 217008 379596 217784 379624
rect 217008 379584 217014 379596
rect 217778 379584 217784 379596
rect 217836 379584 217842 379636
rect 218054 379584 218060 379636
rect 218112 379624 218118 379636
rect 256970 379624 256976 379636
rect 218112 379596 256976 379624
rect 218112 379584 218118 379596
rect 256970 379584 256976 379596
rect 257028 379584 257034 379636
rect 375006 379584 375012 379636
rect 375064 379624 375070 379636
rect 381170 379624 381176 379636
rect 375064 379596 381176 379624
rect 375064 379584 375070 379596
rect 381170 379584 381176 379596
rect 381228 379624 381234 379636
rect 426434 379624 426440 379636
rect 381228 379596 426440 379624
rect 381228 379584 381234 379596
rect 426434 379584 426440 379596
rect 426492 379584 426498 379636
rect 212534 379516 212540 379568
rect 212592 379556 212598 379568
rect 258074 379556 258080 379568
rect 212592 379528 258080 379556
rect 212592 379516 212598 379528
rect 258074 379516 258080 379528
rect 258132 379516 258138 379568
rect 376570 379516 376576 379568
rect 376628 379556 376634 379568
rect 434346 379556 434352 379568
rect 376628 379528 434352 379556
rect 376628 379516 376634 379528
rect 434346 379516 434352 379528
rect 434404 379516 434410 379568
rect 87690 379448 87696 379500
rect 87748 379488 87754 379500
rect 209866 379488 209872 379500
rect 87748 379460 209872 379488
rect 87748 379448 87754 379460
rect 209866 379448 209872 379460
rect 209924 379448 209930 379500
rect 211338 379448 211344 379500
rect 211396 379488 211402 379500
rect 213362 379488 213368 379500
rect 211396 379460 213368 379488
rect 211396 379448 211402 379460
rect 213362 379448 213368 379460
rect 213420 379448 213426 379500
rect 214098 379448 214104 379500
rect 214156 379488 214162 379500
rect 219802 379488 219808 379500
rect 214156 379460 219808 379488
rect 214156 379448 214162 379460
rect 219802 379448 219808 379460
rect 219860 379488 219866 379500
rect 273254 379488 273260 379500
rect 219860 379460 273260 379488
rect 219860 379448 219866 379460
rect 273254 379448 273260 379460
rect 273312 379448 273318 379500
rect 274634 379448 274640 379500
rect 274692 379488 274698 379500
rect 323302 379488 323308 379500
rect 274692 379460 323308 379488
rect 274692 379448 274698 379460
rect 323302 379448 323308 379460
rect 323360 379448 323366 379500
rect 325970 379448 325976 379500
rect 326028 379488 326034 379500
rect 356606 379488 356612 379500
rect 326028 379460 356612 379488
rect 326028 379448 326034 379460
rect 356606 379448 356612 379460
rect 356664 379448 356670 379500
rect 364794 379448 364800 379500
rect 364852 379488 364858 379500
rect 439038 379488 439044 379500
rect 364852 379460 439044 379488
rect 364852 379448 364858 379460
rect 439038 379448 439044 379460
rect 439096 379448 439102 379500
rect 59630 379380 59636 379432
rect 59688 379420 59694 379432
rect 93486 379420 93492 379432
rect 59688 379392 93492 379420
rect 59688 379380 59694 379392
rect 93486 379380 93492 379392
rect 93544 379380 93550 379432
rect 202690 379380 202696 379432
rect 202748 379420 202754 379432
rect 206922 379420 206928 379432
rect 202748 379392 206928 379420
rect 202748 379380 202754 379392
rect 206922 379380 206928 379392
rect 206980 379420 206986 379432
rect 268654 379420 268660 379432
rect 206980 379392 268660 379420
rect 206980 379380 206986 379392
rect 268654 379380 268660 379392
rect 268712 379380 268718 379432
rect 309042 379380 309048 379432
rect 309100 379420 309106 379432
rect 315758 379420 315764 379432
rect 309100 379392 315764 379420
rect 309100 379380 309106 379392
rect 315758 379380 315764 379392
rect 315816 379380 315822 379432
rect 375374 379380 375380 379432
rect 375432 379420 375438 379432
rect 435726 379420 435732 379432
rect 375432 379392 435732 379420
rect 375432 379380 375438 379392
rect 435726 379380 435732 379392
rect 435784 379380 435790 379432
rect 48866 379312 48872 379364
rect 48924 379352 48930 379364
rect 88334 379352 88340 379364
rect 48924 379324 88340 379352
rect 48924 379312 48930 379324
rect 88334 379312 88340 379324
rect 88392 379312 88398 379364
rect 88794 379312 88800 379364
rect 88852 379352 88858 379364
rect 209774 379352 209780 379364
rect 88852 379324 209780 379352
rect 88852 379312 88858 379324
rect 209774 379312 209780 379324
rect 209832 379352 209838 379364
rect 219618 379352 219624 379364
rect 209832 379324 219624 379352
rect 209832 379312 209838 379324
rect 219618 379312 219624 379324
rect 219676 379312 219682 379364
rect 219710 379312 219716 379364
rect 219768 379352 219774 379364
rect 220262 379352 220268 379364
rect 219768 379324 220268 379352
rect 219768 379312 219774 379324
rect 220262 379312 220268 379324
rect 220320 379352 220326 379364
rect 271046 379352 271052 379364
rect 220320 379324 271052 379352
rect 220320 379312 220326 379324
rect 271046 379312 271052 379324
rect 271104 379312 271110 379364
rect 301498 379312 301504 379364
rect 301556 379352 301562 379364
rect 313366 379352 313372 379364
rect 301556 379324 313372 379352
rect 301556 379312 301562 379324
rect 313366 379312 313372 379324
rect 313424 379312 313430 379364
rect 371142 379312 371148 379364
rect 371200 379352 371206 379364
rect 375190 379352 375196 379364
rect 371200 379324 375196 379352
rect 371200 379312 371206 379324
rect 375190 379312 375196 379324
rect 375248 379312 375254 379364
rect 375282 379312 375288 379364
rect 375340 379352 375346 379364
rect 408310 379352 408316 379364
rect 375340 379324 408316 379352
rect 375340 379312 375346 379324
rect 408310 379312 408316 379324
rect 408368 379312 408374 379364
rect 55950 379244 55956 379296
rect 56008 379284 56014 379296
rect 90634 379284 90640 379296
rect 56008 379256 90640 379284
rect 56008 379244 56014 379256
rect 90634 379244 90640 379256
rect 90692 379244 90698 379296
rect 91370 379244 91376 379296
rect 91428 379284 91434 379296
rect 211246 379284 211252 379296
rect 91428 379256 211252 379284
rect 91428 379244 91434 379256
rect 211246 379244 211252 379256
rect 211304 379244 211310 379296
rect 212534 379244 212540 379296
rect 212592 379284 212598 379296
rect 212902 379284 212908 379296
rect 212592 379256 212908 379284
rect 212592 379244 212598 379256
rect 212902 379244 212908 379256
rect 212960 379244 212966 379296
rect 213362 379244 213368 379296
rect 213420 379284 213426 379296
rect 253382 379284 253388 379296
rect 213420 379256 253388 379284
rect 213420 379244 213426 379256
rect 253382 379244 253388 379256
rect 253440 379244 253446 379296
rect 293954 379244 293960 379296
rect 294012 379284 294018 379296
rect 310974 379284 310980 379296
rect 294012 379256 310980 379284
rect 294012 379244 294018 379256
rect 310974 379244 310980 379256
rect 311032 379244 311038 379296
rect 92382 379176 92388 379228
rect 92440 379216 92446 379228
rect 201402 379216 201408 379228
rect 92440 379188 201408 379216
rect 92440 379176 92446 379188
rect 201402 379176 201408 379188
rect 201460 379176 201466 379228
rect 209866 379176 209872 379228
rect 209924 379216 209930 379228
rect 219802 379216 219808 379228
rect 209924 379188 219808 379216
rect 209924 379176 209930 379188
rect 219802 379176 219808 379188
rect 219860 379216 219866 379228
rect 220722 379216 220728 379228
rect 219860 379188 220728 379216
rect 219860 379176 219866 379188
rect 220722 379176 220728 379188
rect 220780 379176 220786 379228
rect 46198 379108 46204 379160
rect 46256 379148 46262 379160
rect 108206 379148 108212 379160
rect 46256 379120 108212 379148
rect 46256 379108 46262 379120
rect 108206 379108 108212 379120
rect 108264 379108 108270 379160
rect 114462 379108 114468 379160
rect 114520 379148 114526 379160
rect 219894 379148 219900 379160
rect 114520 379120 219900 379148
rect 114520 379108 114526 379120
rect 219894 379108 219900 379120
rect 219952 379148 219958 379160
rect 220906 379148 220912 379160
rect 219952 379120 220912 379148
rect 219952 379108 219958 379120
rect 220906 379108 220912 379120
rect 220964 379108 220970 379160
rect 43990 379040 43996 379092
rect 44048 379080 44054 379092
rect 105262 379080 105268 379092
rect 44048 379052 105268 379080
rect 44048 379040 44054 379052
rect 105262 379040 105268 379052
rect 105320 379040 105326 379092
rect 117130 379040 117136 379092
rect 117188 379080 117194 379092
rect 117188 379052 205634 379080
rect 117188 379040 117194 379052
rect 44910 378972 44916 379024
rect 44968 379012 44974 379024
rect 46198 379012 46204 379024
rect 44968 378984 46204 379012
rect 44968 378972 44974 378984
rect 46198 378972 46204 378984
rect 46256 378972 46262 379024
rect 50154 378972 50160 379024
rect 50212 379012 50218 379024
rect 98454 379012 98460 379024
rect 50212 378984 98460 379012
rect 50212 378972 50218 378984
rect 98454 378972 98460 378984
rect 98512 378972 98518 379024
rect 112622 378972 112628 379024
rect 112680 379012 112686 379024
rect 205606 379012 205634 379052
rect 211246 379040 211252 379092
rect 211304 379080 211310 379092
rect 221182 379080 221188 379092
rect 211304 379052 221188 379080
rect 211304 379040 211310 379052
rect 221182 379040 221188 379052
rect 221240 379080 221246 379092
rect 222010 379080 222016 379092
rect 221240 379052 222016 379080
rect 221240 379040 221246 379052
rect 222010 379040 222016 379052
rect 222068 379040 222074 379092
rect 209682 379012 209688 379024
rect 112680 378984 200114 379012
rect 205606 378984 209688 379012
rect 112680 378972 112686 378984
rect 57146 378904 57152 378956
rect 57204 378944 57210 378956
rect 103514 378944 103520 378956
rect 57204 378916 103520 378944
rect 57204 378904 57210 378916
rect 103514 378904 103520 378916
rect 103572 378904 103578 378956
rect 55766 378836 55772 378888
rect 55824 378876 55830 378888
rect 101030 378876 101036 378888
rect 55824 378848 101036 378876
rect 55824 378836 55830 378848
rect 101030 378836 101036 378848
rect 101088 378836 101094 378888
rect 44818 378768 44824 378820
rect 44876 378808 44882 378820
rect 48866 378808 48872 378820
rect 44876 378780 48872 378808
rect 44876 378768 44882 378780
rect 48866 378768 48872 378780
rect 48924 378768 48930 378820
rect 90082 378768 90088 378820
rect 90140 378808 90146 378820
rect 199010 378808 199016 378820
rect 90140 378780 199016 378808
rect 90140 378768 90146 378780
rect 199010 378768 199016 378780
rect 199068 378768 199074 378820
rect 200086 378808 200114 378984
rect 209682 378972 209688 378984
rect 209740 379012 209746 379024
rect 220998 379012 221004 379024
rect 209740 378984 221004 379012
rect 209740 378972 209746 378984
rect 220998 378972 221004 378984
rect 221056 379012 221062 379024
rect 221056 378984 229094 379012
rect 221056 378972 221062 378984
rect 208946 378904 208952 378956
rect 209004 378944 209010 378956
rect 219710 378944 219716 378956
rect 209004 378916 219716 378944
rect 209004 378904 209010 378916
rect 219710 378904 219716 378916
rect 219768 378904 219774 378956
rect 201402 378836 201408 378888
rect 201460 378876 201466 378888
rect 220814 378876 220820 378888
rect 201460 378848 220820 378876
rect 201460 378836 201466 378848
rect 220814 378836 220820 378848
rect 220872 378876 220878 378888
rect 222102 378876 222108 378888
rect 220872 378848 222108 378876
rect 220872 378836 220878 378848
rect 222102 378836 222108 378848
rect 222160 378836 222166 378888
rect 229066 378876 229094 378984
rect 372430 378972 372436 379024
rect 372488 379012 372494 379024
rect 380986 379012 380992 379024
rect 372488 378984 380992 379012
rect 372488 378972 372494 378984
rect 380986 378972 380992 378984
rect 381044 378972 381050 379024
rect 379790 378904 379796 378956
rect 379848 378944 379854 378956
rect 397086 378944 397092 378956
rect 379848 378916 397092 378944
rect 379848 378904 379854 378916
rect 397086 378904 397092 378916
rect 397144 378904 397150 378956
rect 276934 378876 276940 378888
rect 229066 378848 276940 378876
rect 276934 378836 276940 378848
rect 276992 378836 276998 378888
rect 361482 378836 361488 378888
rect 361540 378876 361546 378888
rect 380894 378876 380900 378888
rect 361540 378848 380900 378876
rect 361540 378836 361546 378848
rect 380894 378836 380900 378848
rect 380952 378836 380958 378888
rect 205450 378808 205456 378820
rect 200086 378780 205456 378808
rect 205450 378768 205456 378780
rect 205508 378808 205514 378820
rect 210326 378808 210332 378820
rect 205508 378780 210332 378808
rect 205508 378768 205514 378780
rect 210326 378768 210332 378780
rect 210384 378768 210390 378820
rect 212534 378768 212540 378820
rect 212592 378808 212598 378820
rect 213454 378808 213460 378820
rect 212592 378780 213460 378808
rect 212592 378768 212598 378780
rect 213454 378768 213460 378780
rect 213512 378808 213518 378820
rect 219158 378808 219164 378820
rect 213512 378780 219164 378808
rect 213512 378768 213518 378780
rect 219158 378768 219164 378780
rect 219216 378808 219222 378820
rect 245378 378808 245384 378820
rect 219216 378780 245384 378808
rect 219216 378768 219222 378780
rect 245378 378768 245384 378780
rect 245436 378768 245442 378820
rect 359550 378768 359556 378820
rect 359608 378808 359614 378820
rect 375466 378808 375472 378820
rect 359608 378780 375472 378808
rect 359608 378768 359614 378780
rect 375466 378768 375472 378780
rect 375524 378768 375530 378820
rect 379514 378768 379520 378820
rect 379572 378808 379578 378820
rect 379974 378808 379980 378820
rect 379572 378780 379980 378808
rect 379572 378768 379578 378780
rect 379974 378768 379980 378780
rect 380032 378808 380038 378820
rect 403618 378808 403624 378820
rect 380032 378780 403624 378808
rect 380032 378768 380038 378780
rect 403618 378768 403624 378780
rect 403676 378768 403682 378820
rect 47854 378700 47860 378752
rect 47912 378740 47918 378752
rect 96062 378740 96068 378752
rect 47912 378712 96068 378740
rect 47912 378700 47918 378712
rect 96062 378700 96068 378712
rect 96120 378700 96126 378752
rect 219710 378700 219716 378752
rect 219768 378740 219774 378752
rect 219894 378740 219900 378752
rect 219768 378712 219900 378740
rect 219768 378700 219774 378712
rect 219894 378700 219900 378712
rect 219952 378740 219958 378752
rect 246022 378740 246028 378752
rect 219952 378712 246028 378740
rect 219952 378700 219958 378712
rect 246022 378700 246028 378712
rect 246080 378700 246086 378752
rect 375190 378700 375196 378752
rect 375248 378740 375254 378752
rect 375248 378712 383654 378740
rect 375248 378700 375254 378712
rect 86586 378632 86592 378684
rect 86644 378672 86650 378684
rect 208946 378672 208952 378684
rect 86644 378644 208952 378672
rect 86644 378632 86650 378644
rect 208946 378632 208952 378644
rect 209004 378632 209010 378684
rect 220722 378632 220728 378684
rect 220780 378672 220786 378684
rect 247494 378672 247500 378684
rect 220780 378644 247500 378672
rect 220780 378632 220786 378644
rect 247494 378632 247500 378644
rect 247552 378632 247558 378684
rect 383626 378672 383654 378712
rect 396074 378672 396080 378684
rect 383626 378644 396080 378672
rect 396074 378632 396080 378644
rect 396132 378632 396138 378684
rect 199010 378564 199016 378616
rect 199068 378604 199074 378616
rect 221274 378604 221280 378616
rect 199068 378576 221280 378604
rect 199068 378564 199074 378576
rect 221274 378564 221280 378576
rect 221332 378604 221338 378616
rect 250070 378604 250076 378616
rect 221332 378576 250076 378604
rect 221332 378564 221338 378576
rect 250070 378564 250076 378576
rect 250128 378564 250134 378616
rect 379330 378564 379336 378616
rect 379388 378604 379394 378616
rect 379514 378604 379520 378616
rect 379388 378576 379520 378604
rect 379388 378564 379394 378576
rect 379514 378564 379520 378576
rect 379572 378604 379578 378616
rect 405826 378604 405832 378616
rect 379572 378576 405832 378604
rect 379572 378564 379578 378576
rect 405826 378564 405832 378576
rect 405884 378564 405890 378616
rect 219618 378496 219624 378548
rect 219676 378536 219682 378548
rect 248598 378536 248604 378548
rect 219676 378508 248604 378536
rect 219676 378496 219682 378508
rect 248598 378496 248604 378508
rect 248656 378496 248662 378548
rect 380986 378496 380992 378548
rect 381044 378536 381050 378548
rect 412358 378536 412364 378548
rect 381044 378508 412364 378536
rect 381044 378496 381050 378508
rect 412358 378496 412364 378508
rect 412416 378496 412422 378548
rect 108850 378428 108856 378480
rect 108908 378468 108914 378480
rect 202690 378468 202696 378480
rect 108908 378440 202696 378468
rect 108908 378428 108914 378440
rect 202690 378428 202696 378440
rect 202748 378428 202754 378480
rect 210234 378428 210240 378480
rect 210292 378468 210298 378480
rect 211338 378468 211344 378480
rect 210292 378440 211344 378468
rect 210292 378428 210298 378440
rect 211338 378428 211344 378440
rect 211396 378428 211402 378480
rect 222010 378428 222016 378480
rect 222068 378468 222074 378480
rect 251174 378468 251180 378480
rect 222068 378440 251180 378468
rect 222068 378428 222074 378440
rect 251174 378428 251180 378440
rect 251232 378428 251238 378480
rect 380894 378428 380900 378480
rect 380952 378468 380958 378480
rect 411254 378468 411260 378480
rect 380952 378440 411260 378468
rect 380952 378428 380958 378440
rect 411254 378428 411260 378440
rect 411312 378428 411318 378480
rect 113450 378360 113456 378412
rect 113508 378400 113514 378412
rect 214098 378400 214104 378412
rect 113508 378372 214104 378400
rect 113508 378360 113514 378372
rect 214098 378360 214104 378372
rect 214156 378360 214162 378412
rect 222102 378360 222108 378412
rect 222160 378400 222166 378412
rect 252278 378400 252284 378412
rect 222160 378372 252284 378400
rect 222160 378360 222166 378372
rect 252278 378360 252284 378372
rect 252336 378360 252342 378412
rect 343450 378360 343456 378412
rect 343508 378400 343514 378412
rect 357526 378400 357532 378412
rect 343508 378372 357532 378400
rect 343508 378360 343514 378372
rect 357526 378360 357532 378372
rect 357584 378400 357590 378412
rect 358630 378400 358636 378412
rect 357584 378372 358636 378400
rect 357584 378360 357590 378372
rect 358630 378360 358636 378372
rect 358688 378360 358694 378412
rect 375466 378360 375472 378412
rect 375524 378400 375530 378412
rect 376386 378400 376392 378412
rect 375524 378372 376392 378400
rect 375524 378360 375530 378372
rect 376386 378360 376392 378372
rect 376444 378400 376450 378412
rect 407574 378400 407580 378412
rect 376444 378372 407580 378400
rect 376444 378360 376450 378372
rect 407574 378360 407580 378372
rect 407632 378360 407638 378412
rect 111242 378292 111248 378344
rect 111300 378332 111306 378344
rect 213362 378332 213368 378344
rect 111300 378304 213368 378332
rect 111300 378292 111306 378304
rect 213362 378292 213368 378304
rect 213420 378332 213426 378344
rect 220262 378332 220268 378344
rect 213420 378304 220268 378332
rect 213420 378292 213426 378304
rect 220262 378292 220268 378304
rect 220320 378292 220326 378344
rect 220906 378292 220912 378344
rect 220964 378332 220970 378344
rect 274174 378332 274180 378344
rect 220964 378304 274180 378332
rect 220964 378292 220970 378304
rect 274174 378292 274180 378304
rect 274232 378292 274238 378344
rect 274266 378292 274272 378344
rect 274324 378332 274330 378344
rect 302786 378332 302792 378344
rect 274324 378304 302792 378332
rect 274324 378292 274330 378304
rect 302786 378292 302792 378304
rect 302844 378292 302850 378344
rect 342254 378292 342260 378344
rect 342312 378332 342318 378344
rect 343174 378332 343180 378344
rect 342312 378304 343180 378332
rect 342312 378292 342318 378304
rect 343174 378292 343180 378304
rect 343232 378332 343238 378344
rect 359366 378332 359372 378344
rect 343232 378304 359372 378332
rect 343232 378292 343238 378304
rect 359366 378292 359372 378304
rect 359424 378332 359430 378344
rect 359424 378304 364334 378332
rect 359424 378292 359430 378304
rect 48866 378224 48872 378276
rect 48924 378264 48930 378276
rect 81434 378264 81440 378276
rect 48924 378236 81440 378264
rect 48924 378224 48930 378236
rect 81434 378224 81440 378236
rect 81492 378224 81498 378276
rect 93394 378224 93400 378276
rect 93452 378264 93458 378276
rect 210234 378264 210240 378276
rect 93452 378236 210240 378264
rect 93452 378224 93458 378236
rect 210234 378224 210240 378236
rect 210292 378224 210298 378276
rect 210326 378224 210332 378276
rect 210384 378264 210390 378276
rect 272058 378264 272064 378276
rect 210384 378236 272064 378264
rect 210384 378224 210390 378236
rect 272058 378224 272064 378236
rect 272116 378224 272122 378276
rect 277854 378224 277860 378276
rect 277912 378264 277918 378276
rect 357434 378264 357440 378276
rect 277912 378236 357440 378264
rect 277912 378224 277918 378236
rect 357434 378224 357440 378236
rect 357492 378224 357498 378276
rect 364306 378264 364334 378304
rect 377122 378292 377128 378344
rect 377180 378332 377186 378344
rect 379422 378332 379428 378344
rect 377180 378304 379428 378332
rect 377180 378292 377186 378304
rect 379422 378292 379428 378304
rect 379480 378332 379486 378344
rect 426618 378332 426624 378344
rect 379480 378304 426624 378332
rect 379480 378292 379486 378304
rect 426618 378292 426624 378304
rect 426676 378292 426682 378344
rect 439038 378292 439044 378344
rect 439096 378332 439102 378344
rect 516594 378332 516600 378344
rect 439096 378304 516600 378332
rect 439096 378292 439102 378304
rect 516594 378292 516600 378304
rect 516652 378292 516658 378344
rect 503070 378264 503076 378276
rect 364306 378236 503076 378264
rect 503070 378224 503076 378236
rect 503128 378264 503134 378276
rect 517606 378264 517612 378276
rect 503128 378236 517612 378264
rect 503128 378224 503134 378236
rect 517606 378224 517612 378236
rect 517664 378264 517670 378276
rect 580258 378264 580264 378276
rect 517664 378236 580264 378264
rect 517664 378224 517670 378236
rect 580258 378224 580264 378236
rect 580316 378224 580322 378276
rect 46198 378156 46204 378208
rect 46256 378196 46262 378208
rect 80422 378196 80428 378208
rect 46256 378168 80428 378196
rect 46256 378156 46262 378168
rect 80422 378156 80428 378168
rect 80480 378156 80486 378208
rect 85482 378156 85488 378208
rect 85540 378196 85546 378208
rect 212534 378196 212540 378208
rect 85540 378168 212540 378196
rect 85540 378156 85546 378168
rect 212534 378156 212540 378168
rect 212592 378156 212598 378208
rect 274634 378156 274640 378208
rect 274692 378196 274698 378208
rect 275646 378196 275652 378208
rect 274692 378168 275652 378196
rect 274692 378156 274698 378168
rect 275646 378156 275652 378168
rect 275704 378196 275710 378208
rect 356606 378196 356612 378208
rect 275704 378168 356612 378196
rect 275704 378156 275710 378168
rect 356606 378156 356612 378168
rect 356664 378156 356670 378208
rect 358630 378156 358636 378208
rect 358688 378196 358694 378208
rect 503530 378196 503536 378208
rect 358688 378168 503536 378196
rect 358688 378156 358694 378168
rect 503530 378156 503536 378168
rect 503588 378196 503594 378208
rect 517698 378196 517704 378208
rect 503588 378168 517704 378196
rect 503588 378156 503594 378168
rect 517698 378156 517704 378168
rect 517756 378196 517762 378208
rect 580166 378196 580172 378208
rect 517756 378168 580172 378196
rect 517756 378156 517762 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 43254 378088 43260 378140
rect 43312 378128 43318 378140
rect 199102 378128 199108 378140
rect 43312 378100 199108 378128
rect 43312 378088 43318 378100
rect 199102 378088 199108 378100
rect 199160 378128 199166 378140
rect 199838 378128 199844 378140
rect 199160 378100 199844 378128
rect 199160 378088 199166 378100
rect 199838 378088 199844 378100
rect 199896 378088 199902 378140
rect 201494 378088 201500 378140
rect 201552 378128 201558 378140
rect 317414 378128 317420 378140
rect 201552 378100 317420 378128
rect 201552 378088 201558 378100
rect 317414 378088 317420 378100
rect 317472 378088 317478 378140
rect 357066 378088 357072 378140
rect 357124 378128 357130 378140
rect 474826 378128 474832 378140
rect 357124 378100 474832 378128
rect 357124 378088 357130 378100
rect 474826 378088 474832 378100
rect 474884 378088 474890 378140
rect 54386 378020 54392 378072
rect 54444 378060 54450 378072
rect 183186 378060 183192 378072
rect 54444 378032 183192 378060
rect 54444 378020 54450 378032
rect 183186 378020 183192 378032
rect 183244 378060 183250 378072
rect 197998 378060 198004 378072
rect 183244 378032 198004 378060
rect 183244 378020 183250 378032
rect 197998 378020 198004 378032
rect 198056 378020 198062 378072
rect 198826 378020 198832 378072
rect 198884 378060 198890 378072
rect 300854 378060 300860 378072
rect 198884 378032 300860 378060
rect 198884 378020 198890 378032
rect 300854 378020 300860 378032
rect 300912 378020 300918 378072
rect 358722 378020 358728 378072
rect 358780 378060 358786 378072
rect 460934 378060 460940 378072
rect 358780 378032 460940 378060
rect 358780 378020 358786 378032
rect 460934 378020 460940 378032
rect 460992 378020 460998 378072
rect 54294 377952 54300 378004
rect 54352 377992 54358 378004
rect 182266 377992 182272 378004
rect 54352 377964 182272 377992
rect 54352 377952 54358 377964
rect 182266 377952 182272 377964
rect 182324 377952 182330 378004
rect 197446 377952 197452 378004
rect 197504 377992 197510 378004
rect 298462 377992 298468 378004
rect 197504 377964 298468 377992
rect 197504 377952 197510 377964
rect 298462 377952 298468 377964
rect 298520 377952 298526 378004
rect 374362 377952 374368 378004
rect 374420 377992 374426 378004
rect 458358 377992 458364 378004
rect 374420 377964 458364 377992
rect 374420 377952 374426 377964
rect 458358 377952 458364 377964
rect 458416 377952 458422 378004
rect 105538 377884 105544 377936
rect 105596 377924 105602 377936
rect 215386 377924 215392 377936
rect 105596 377896 215392 377924
rect 105596 377884 105602 377896
rect 215386 377884 215392 377896
rect 215444 377924 215450 377936
rect 215754 377924 215760 377936
rect 215444 377896 215760 377924
rect 215444 377884 215450 377896
rect 215754 377884 215760 377896
rect 215812 377884 215818 377936
rect 217502 377884 217508 377936
rect 217560 377924 217566 377936
rect 305822 377924 305828 377936
rect 217560 377896 305828 377924
rect 217560 377884 217566 377896
rect 305822 377884 305828 377896
rect 305880 377884 305886 377936
rect 370314 377884 370320 377936
rect 370372 377924 370378 377936
rect 452746 377924 452752 377936
rect 370372 377896 452752 377924
rect 370372 377884 370378 377896
rect 452746 377884 452752 377896
rect 452804 377884 452810 377936
rect 150986 377816 150992 377868
rect 151044 377856 151050 377868
rect 198090 377856 198096 377868
rect 151044 377828 198096 377856
rect 151044 377816 151050 377828
rect 198090 377816 198096 377828
rect 198148 377816 198154 377868
rect 198274 377816 198280 377868
rect 198332 377856 198338 377868
rect 295886 377856 295892 377868
rect 198332 377828 295892 377856
rect 198332 377816 198338 377828
rect 295886 377816 295892 377828
rect 295944 377816 295950 377868
rect 365438 377816 365444 377868
rect 365496 377856 365502 377868
rect 447502 377856 447508 377868
rect 365496 377828 447508 377856
rect 365496 377816 365502 377828
rect 447502 377816 447508 377828
rect 447560 377816 447566 377868
rect 148594 377748 148600 377800
rect 148652 377788 148658 377800
rect 197262 377788 197268 377800
rect 148652 377760 197268 377788
rect 148652 377748 148658 377760
rect 197262 377748 197268 377760
rect 197320 377748 197326 377800
rect 197538 377748 197544 377800
rect 197596 377788 197602 377800
rect 292666 377788 292672 377800
rect 197596 377760 292672 377788
rect 197596 377748 197602 377760
rect 292666 377748 292672 377760
rect 292724 377748 292730 377800
rect 373718 377748 373724 377800
rect 373776 377788 373782 377800
rect 455598 377788 455604 377800
rect 373776 377760 455604 377788
rect 373776 377748 373782 377760
rect 455598 377748 455604 377760
rect 455656 377748 455662 377800
rect 196710 377680 196716 377732
rect 196768 377720 196774 377732
rect 290918 377720 290924 377732
rect 196768 377692 290924 377720
rect 196768 377680 196774 377692
rect 290918 377680 290924 377692
rect 290976 377680 290982 377732
rect 450998 377720 451004 377732
rect 371804 377692 451004 377720
rect 196802 377612 196808 377664
rect 196860 377652 196866 377664
rect 287698 377652 287704 377664
rect 196860 377624 287704 377652
rect 196860 377612 196866 377624
rect 287698 377612 287704 377624
rect 287756 377612 287762 377664
rect 359458 377612 359464 377664
rect 359516 377652 359522 377664
rect 369854 377652 369860 377664
rect 359516 377624 369860 377652
rect 359516 377612 359522 377624
rect 369854 377612 369860 377624
rect 369912 377612 369918 377664
rect 196618 377544 196624 377596
rect 196676 377584 196682 377596
rect 285950 377584 285956 377596
rect 196676 377556 285956 377584
rect 196676 377544 196682 377556
rect 285950 377544 285956 377556
rect 286008 377544 286014 377596
rect 368382 377544 368388 377596
rect 368440 377584 368446 377596
rect 371804 377584 371832 377692
rect 450998 377680 451004 377692
rect 451056 377680 451062 377732
rect 423398 377652 423404 377664
rect 368440 377556 371832 377584
rect 371988 377624 423404 377652
rect 368440 377544 368446 377556
rect 98270 377476 98276 377528
rect 98328 377516 98334 377528
rect 208946 377516 208952 377528
rect 98328 377488 208952 377516
rect 98328 377476 98334 377488
rect 208946 377476 208952 377488
rect 209004 377516 209010 377528
rect 212902 377516 212908 377528
rect 209004 377488 212908 377516
rect 209004 377476 209010 377488
rect 212902 377476 212908 377488
rect 212960 377476 212966 377528
rect 215754 377476 215760 377528
rect 215812 377516 215818 377528
rect 219342 377516 219348 377528
rect 215812 377488 219348 377516
rect 215812 377476 215818 377488
rect 219342 377476 219348 377488
rect 219400 377516 219406 377528
rect 237374 377516 237380 377528
rect 219400 377488 237380 377516
rect 219400 377476 219406 377488
rect 237374 377476 237380 377488
rect 237432 377476 237438 377528
rect 369854 377476 369860 377528
rect 369912 377516 369918 377528
rect 371988 377516 372016 377624
rect 423398 377612 423404 377624
rect 423456 377612 423462 377664
rect 372798 377544 372804 377596
rect 372856 377584 372862 377596
rect 413094 377584 413100 377596
rect 372856 377556 413100 377584
rect 372856 377544 372862 377556
rect 413094 377544 413100 377556
rect 413152 377544 413158 377596
rect 369912 377488 372016 377516
rect 369912 377476 369918 377488
rect 379882 377476 379888 377528
rect 379940 377516 379946 377528
rect 414566 377516 414572 377528
rect 379940 377488 414572 377516
rect 379940 377476 379946 377488
rect 414566 377476 414572 377488
rect 414624 377476 414630 377528
rect 199378 377408 199384 377460
rect 199436 377448 199442 377460
rect 280706 377448 280712 377460
rect 199436 377420 280712 377448
rect 199436 377408 199442 377420
rect 280706 377408 280712 377420
rect 280764 377408 280770 377460
rect 367002 377408 367008 377460
rect 367060 377448 367066 377460
rect 375282 377448 375288 377460
rect 367060 377420 375288 377448
rect 367060 377408 367066 377420
rect 375282 377408 375288 377420
rect 375340 377408 375346 377460
rect 415762 377448 415768 377460
rect 379486 377420 415768 377448
rect 197078 377340 197084 377392
rect 197136 377380 197142 377392
rect 278038 377380 278044 377392
rect 197136 377352 278044 377380
rect 197136 377340 197142 377352
rect 278038 377340 278044 377352
rect 278096 377340 278102 377392
rect 379486 377380 379514 377420
rect 415762 377408 415768 377420
rect 415820 377408 415826 377460
rect 410058 377380 410064 377392
rect 377232 377352 379514 377380
rect 379900 377352 410064 377380
rect 198734 377272 198740 377324
rect 198792 377312 198798 377324
rect 274266 377312 274272 377324
rect 198792 377284 274272 377312
rect 198792 377272 198798 377284
rect 274266 377272 274272 377284
rect 274324 377272 274330 377324
rect 375282 377272 375288 377324
rect 375340 377312 375346 377324
rect 377232 377312 377260 377352
rect 375340 377284 377260 377312
rect 375340 377272 375346 377284
rect 377306 377272 377312 377324
rect 377364 377312 377370 377324
rect 379900 377312 379928 377352
rect 410058 377340 410064 377352
rect 410116 377340 410122 377392
rect 402974 377312 402980 377324
rect 377364 377284 379928 377312
rect 383626 377284 402980 377312
rect 377364 377272 377370 377284
rect 153562 377204 153568 377256
rect 153620 377244 153626 377256
rect 200390 377244 200396 377256
rect 153620 377216 200396 377244
rect 153620 377204 153626 377216
rect 200390 377204 200396 377216
rect 200448 377204 200454 377256
rect 373902 377204 373908 377256
rect 373960 377244 373966 377256
rect 375926 377244 375932 377256
rect 373960 377216 375932 377244
rect 373960 377204 373966 377216
rect 375926 377204 375932 377216
rect 375984 377244 375990 377256
rect 383626 377244 383654 377284
rect 402974 377272 402980 377284
rect 403032 377272 403038 377324
rect 375984 377216 383654 377244
rect 375984 377204 375990 377216
rect 141050 377136 141056 377188
rect 141108 377176 141114 377188
rect 200482 377176 200488 377188
rect 141108 377148 200488 377176
rect 141108 377136 141114 377148
rect 200482 377136 200488 377148
rect 200540 377136 200546 377188
rect 374454 377136 374460 377188
rect 374512 377176 374518 377188
rect 379882 377176 379888 377188
rect 374512 377148 379888 377176
rect 374512 377136 374518 377148
rect 379882 377136 379888 377148
rect 379940 377136 379946 377188
rect 42150 377068 42156 377120
rect 42208 377108 42214 377120
rect 199470 377108 199476 377120
rect 42208 377080 199476 377108
rect 42208 377068 42214 377080
rect 199470 377068 199476 377080
rect 199528 377068 199534 377120
rect 380894 376932 380900 376984
rect 380952 376972 380958 376984
rect 381170 376972 381176 376984
rect 380952 376944 381176 376972
rect 380952 376932 380958 376944
rect 381170 376932 381176 376944
rect 381228 376932 381234 376984
rect 212994 376660 213000 376712
rect 213052 376700 213058 376712
rect 283006 376700 283012 376712
rect 213052 376672 283012 376700
rect 213052 376660 213058 376672
rect 283006 376660 283012 376672
rect 283064 376660 283070 376712
rect 361298 376660 361304 376712
rect 361356 376700 361362 376712
rect 477586 376700 477592 376712
rect 361356 376672 477592 376700
rect 361356 376660 361362 376672
rect 477586 376660 477592 376672
rect 477644 376660 477650 376712
rect 83458 376592 83464 376644
rect 83516 376632 83522 376644
rect 207106 376632 207112 376644
rect 83516 376604 207112 376632
rect 83516 376592 83522 376604
rect 207106 376592 207112 376604
rect 207164 376592 207170 376644
rect 210142 376592 210148 376644
rect 210200 376632 210206 376644
rect 320910 376632 320916 376644
rect 210200 376604 320916 376632
rect 210200 376592 210206 376604
rect 320910 376592 320916 376604
rect 320968 376592 320974 376644
rect 366266 376592 366272 376644
rect 366324 376632 366330 376644
rect 480530 376632 480536 376644
rect 366324 376604 480536 376632
rect 366324 376592 366330 376604
rect 480530 376592 480536 376604
rect 480588 376592 480594 376644
rect 203886 376524 203892 376576
rect 203944 376564 203950 376576
rect 273438 376564 273444 376576
rect 203944 376536 273444 376564
rect 203944 376524 203950 376536
rect 273438 376524 273444 376536
rect 273496 376524 273502 376576
rect 364150 376524 364156 376576
rect 364208 376564 364214 376576
rect 473446 376564 473452 376576
rect 364208 376536 473452 376564
rect 364208 376524 364214 376536
rect 473446 376524 473452 376536
rect 473504 376524 473510 376576
rect 97166 376456 97172 376508
rect 97224 376496 97230 376508
rect 97224 376468 200114 376496
rect 97224 376456 97230 376468
rect 200086 376360 200114 376468
rect 211614 376456 211620 376508
rect 211672 376496 211678 376508
rect 211672 376468 212856 376496
rect 211672 376456 211678 376468
rect 210050 376388 210056 376440
rect 210108 376428 210114 376440
rect 212626 376428 212632 376440
rect 210108 376400 212632 376428
rect 210108 376388 210114 376400
rect 212626 376388 212632 376400
rect 212684 376388 212690 376440
rect 212534 376360 212540 376372
rect 200086 376332 212540 376360
rect 212534 376320 212540 376332
rect 212592 376320 212598 376372
rect 212828 376360 212856 376468
rect 213914 376456 213920 376508
rect 213972 376496 213978 376508
rect 216398 376496 216404 376508
rect 213972 376468 216404 376496
rect 213972 376456 213978 376468
rect 216398 376456 216404 376468
rect 216456 376456 216462 376508
rect 217594 376456 217600 376508
rect 217652 376496 217658 376508
rect 276014 376496 276020 376508
rect 217652 376468 276020 376496
rect 217652 376456 217658 376468
rect 276014 376456 276020 376468
rect 276072 376456 276078 376508
rect 362678 376456 362684 376508
rect 362736 376496 362742 376508
rect 470870 376496 470876 376508
rect 362736 376468 470876 376496
rect 362736 376456 362742 376468
rect 470870 376456 470876 376468
rect 470928 376456 470934 376508
rect 213546 376388 213552 376440
rect 213604 376428 213610 376440
rect 268102 376428 268108 376440
rect 213604 376400 268108 376428
rect 213604 376388 213610 376400
rect 268102 376388 268108 376400
rect 268160 376388 268166 376440
rect 364702 376388 364708 376440
rect 364760 376428 364766 376440
rect 467926 376428 467932 376440
rect 364760 376400 467932 376428
rect 364760 376388 364766 376400
rect 467926 376388 467932 376400
rect 467984 376388 467990 376440
rect 212828 376332 212948 376360
rect 138474 376252 138480 376304
rect 138532 376292 138538 376304
rect 201770 376292 201776 376304
rect 138532 376264 201776 376292
rect 138532 376252 138538 376264
rect 201770 376252 201776 376264
rect 201828 376252 201834 376304
rect 212920 376292 212948 376332
rect 213086 376320 213092 376372
rect 213144 376360 213150 376372
rect 265894 376360 265900 376372
rect 213144 376332 265900 376360
rect 213144 376320 213150 376332
rect 265894 376320 265900 376332
rect 265952 376320 265958 376372
rect 367646 376320 367652 376372
rect 367704 376360 367710 376372
rect 465074 376360 465080 376372
rect 367704 376332 465080 376360
rect 367704 376320 367710 376332
rect 465074 376320 465080 376332
rect 465132 376320 465138 376372
rect 263594 376292 263600 376304
rect 212920 376264 263600 376292
rect 263594 376252 263600 376264
rect 263652 376252 263658 376304
rect 364242 376252 364248 376304
rect 364300 376292 364306 376304
rect 427906 376292 427912 376304
rect 364300 376264 427912 376292
rect 364300 376252 364306 376264
rect 427906 376252 427912 376264
rect 427964 376252 427970 376304
rect 94682 376184 94688 376236
rect 94740 376224 94746 376236
rect 212718 376224 212724 376236
rect 94740 376196 212724 376224
rect 94740 376184 94746 376196
rect 212718 376184 212724 376196
rect 212776 376184 212782 376236
rect 219250 376184 219256 376236
rect 219308 376224 219314 376236
rect 270954 376224 270960 376236
rect 219308 376196 270960 376224
rect 219308 376184 219314 376196
rect 270954 376184 270960 376196
rect 271012 376184 271018 376236
rect 362770 376184 362776 376236
rect 362828 376224 362834 376236
rect 425974 376224 425980 376236
rect 362828 376196 425980 376224
rect 362828 376184 362834 376196
rect 425974 376184 425980 376196
rect 426032 376184 426038 376236
rect 202506 376116 202512 376168
rect 202564 376156 202570 376168
rect 248230 376156 248236 376168
rect 202564 376128 248236 376156
rect 202564 376116 202570 376128
rect 248230 376116 248236 376128
rect 248288 376116 248294 376168
rect 372522 376116 372528 376168
rect 372580 376156 372586 376168
rect 418246 376156 418252 376168
rect 372580 376128 418252 376156
rect 372580 376116 372586 376128
rect 418246 376116 418252 376128
rect 418304 376116 418310 376168
rect 99466 376048 99472 376100
rect 99524 376088 99530 376100
rect 213914 376088 213920 376100
rect 99524 376060 213920 376088
rect 99524 376048 99530 376060
rect 213914 376048 213920 376060
rect 213972 376048 213978 376100
rect 215846 376048 215852 376100
rect 215904 376088 215910 376100
rect 260926 376088 260932 376100
rect 215904 376060 260932 376088
rect 215904 376048 215910 376060
rect 260926 376048 260932 376060
rect 260984 376048 260990 376100
rect 370406 376048 370412 376100
rect 370464 376088 370470 376100
rect 416038 376088 416044 376100
rect 370464 376060 416044 376088
rect 370464 376048 370470 376060
rect 416038 376048 416044 376060
rect 416096 376048 416102 376100
rect 95970 375980 95976 376032
rect 96028 376020 96034 376032
rect 213730 376020 213736 376032
rect 96028 375992 213736 376020
rect 96028 375980 96034 375992
rect 213730 375980 213736 375992
rect 213788 375980 213794 376032
rect 219526 375980 219532 376032
rect 219584 376020 219590 376032
rect 258350 376020 258356 376032
rect 219584 375992 258356 376020
rect 219584 375980 219590 375992
rect 258350 375980 258356 375992
rect 258408 375980 258414 376032
rect 357158 375980 357164 376032
rect 357216 376020 357222 376032
rect 357216 375992 369854 376020
rect 357216 375980 357222 375992
rect 208762 375912 208768 375964
rect 208820 375952 208826 375964
rect 253566 375952 253572 375964
rect 208820 375924 253572 375952
rect 208820 375912 208826 375924
rect 253566 375912 253572 375924
rect 253624 375912 253630 375964
rect 369826 375952 369854 375992
rect 379238 375980 379244 376032
rect 379296 376020 379302 376032
rect 381170 376020 381176 376032
rect 379296 375992 381176 376020
rect 379296 375980 379302 375992
rect 381170 375980 381176 375992
rect 381228 376020 381234 376032
rect 436462 376020 436468 376032
rect 381228 375992 436468 376020
rect 381228 375980 381234 375992
rect 436462 375980 436468 375992
rect 436520 375980 436526 376032
rect 375834 375952 375840 375964
rect 369826 375924 375840 375952
rect 375834 375912 375840 375924
rect 375892 375952 375898 375964
rect 416958 375952 416964 375964
rect 375892 375924 416964 375952
rect 375892 375912 375898 375924
rect 416958 375912 416964 375924
rect 417016 375912 417022 375964
rect 215018 375844 215024 375896
rect 215076 375884 215082 375896
rect 250622 375884 250628 375896
rect 215076 375856 250628 375884
rect 215076 375844 215082 375856
rect 250622 375844 250628 375856
rect 250680 375844 250686 375896
rect 216766 375816 216772 375828
rect 200086 375788 216772 375816
rect 44634 375708 44640 375760
rect 44692 375748 44698 375760
rect 200086 375748 200114 375788
rect 216766 375776 216772 375788
rect 216824 375816 216830 375828
rect 217594 375816 217600 375828
rect 216824 375788 217600 375816
rect 216824 375776 216830 375788
rect 217594 375776 217600 375788
rect 217652 375776 217658 375828
rect 240042 375816 240048 375828
rect 219406 375788 240048 375816
rect 44692 375720 200114 375748
rect 44692 375708 44698 375720
rect 104434 375640 104440 375692
rect 104492 375680 104498 375692
rect 216582 375680 216588 375692
rect 104492 375652 216588 375680
rect 104492 375640 104498 375652
rect 216582 375640 216588 375652
rect 216640 375680 216646 375692
rect 217226 375680 217232 375692
rect 216640 375652 217232 375680
rect 216640 375640 216646 375652
rect 217226 375640 217232 375652
rect 217284 375640 217290 375692
rect 212534 375572 212540 375624
rect 212592 375612 212598 375624
rect 214374 375612 214380 375624
rect 212592 375584 214380 375612
rect 212592 375572 212598 375584
rect 214374 375572 214380 375584
rect 214432 375612 214438 375624
rect 214926 375612 214932 375624
rect 214432 375584 214932 375612
rect 214432 375572 214438 375584
rect 214926 375572 214932 375584
rect 214984 375572 214990 375624
rect 216398 375572 216404 375624
rect 216456 375612 216462 375624
rect 219406 375612 219434 375788
rect 240042 375776 240048 375788
rect 240100 375776 240106 375828
rect 216456 375584 219434 375612
rect 216456 375572 216462 375584
rect 213546 375368 213552 375420
rect 213604 375408 213610 375420
rect 213730 375408 213736 375420
rect 213604 375380 213736 375408
rect 213604 375368 213610 375380
rect 213730 375368 213736 375380
rect 213788 375368 213794 375420
rect 357158 375408 357164 375420
rect 280080 375380 357164 375408
rect 107562 375300 107568 375352
rect 107620 375340 107626 375352
rect 208302 375340 208308 375352
rect 107620 375312 208308 375340
rect 107620 375300 107626 375312
rect 208302 375300 208308 375312
rect 208360 375340 208366 375352
rect 217502 375340 217508 375352
rect 208360 375312 217508 375340
rect 208360 375300 208366 375312
rect 217502 375300 217508 375312
rect 217560 375340 217566 375352
rect 217560 375312 219434 375340
rect 217560 375300 217566 375312
rect 106458 375232 106464 375284
rect 106516 375272 106522 375284
rect 208026 375272 208032 375284
rect 106516 375244 208032 375272
rect 106516 375232 106522 375244
rect 208026 375232 208032 375244
rect 208084 375232 208090 375284
rect 219406 375272 219434 375312
rect 267550 375272 267556 375284
rect 219406 375244 267556 375272
rect 267550 375232 267556 375244
rect 267608 375232 267614 375284
rect 102962 375164 102968 375216
rect 103020 375204 103026 375216
rect 215294 375204 215300 375216
rect 103020 375176 215300 375204
rect 103020 375164 103026 375176
rect 215294 375164 215300 375176
rect 215352 375204 215358 375216
rect 216582 375204 216588 375216
rect 215352 375176 216588 375204
rect 215352 375164 215358 375176
rect 216582 375164 216588 375176
rect 216640 375204 216646 375216
rect 262766 375204 262772 375216
rect 216640 375176 262772 375204
rect 216640 375164 216646 375176
rect 262766 375164 262772 375176
rect 262824 375164 262830 375216
rect 101858 375096 101864 375148
rect 101916 375136 101922 375148
rect 214466 375136 214472 375148
rect 101916 375108 214472 375136
rect 101916 375096 101922 375108
rect 214466 375096 214472 375108
rect 214524 375136 214530 375148
rect 261662 375136 261668 375148
rect 214524 375108 261668 375136
rect 214524 375096 214530 375108
rect 261662 375096 261668 375108
rect 261720 375096 261726 375148
rect 208118 375028 208124 375080
rect 208176 375068 208182 375080
rect 279142 375068 279148 375080
rect 208176 375040 279148 375068
rect 208176 375028 208182 375040
rect 279142 375028 279148 375040
rect 279200 375068 279206 375080
rect 280080 375068 280108 375380
rect 357158 375368 357164 375380
rect 357216 375368 357222 375420
rect 368382 375368 368388 375420
rect 368440 375408 368446 375420
rect 371234 375408 371240 375420
rect 368440 375380 371240 375408
rect 368440 375368 368446 375380
rect 371234 375368 371240 375380
rect 371292 375408 371298 375420
rect 372522 375408 372528 375420
rect 371292 375380 372528 375408
rect 371292 375368 371298 375380
rect 372522 375368 372528 375380
rect 372580 375368 372586 375420
rect 370222 375300 370228 375352
rect 370280 375340 370286 375352
rect 431126 375340 431132 375352
rect 370280 375312 431132 375340
rect 370280 375300 370286 375312
rect 431126 375300 431132 375312
rect 431184 375300 431190 375352
rect 364058 375232 364064 375284
rect 364116 375272 364122 375284
rect 377950 375272 377956 375284
rect 364116 375244 377956 375272
rect 364116 375232 364122 375244
rect 377950 375232 377956 375244
rect 378008 375272 378014 375284
rect 437750 375272 437756 375284
rect 378008 375244 437756 375272
rect 378008 375232 378014 375244
rect 437750 375232 437756 375244
rect 437808 375232 437814 375284
rect 369762 375164 369768 375216
rect 369820 375204 369826 375216
rect 371786 375204 371792 375216
rect 369820 375176 371792 375204
rect 369820 375164 369826 375176
rect 371786 375164 371792 375176
rect 371844 375164 371850 375216
rect 373810 375164 373816 375216
rect 373868 375204 373874 375216
rect 432230 375204 432236 375216
rect 373868 375176 432236 375204
rect 373868 375164 373874 375176
rect 432230 375164 432236 375176
rect 432288 375164 432294 375216
rect 372522 375096 372528 375148
rect 372580 375136 372586 375148
rect 428274 375136 428280 375148
rect 372580 375108 428280 375136
rect 372580 375096 372586 375108
rect 428274 375096 428280 375108
rect 428332 375096 428338 375148
rect 279200 375040 280108 375068
rect 279200 375028 279206 375040
rect 364886 375028 364892 375080
rect 364944 375068 364950 375080
rect 378134 375068 378140 375080
rect 364944 375040 378140 375068
rect 364944 375028 364950 375040
rect 378134 375028 378140 375040
rect 378192 375028 378198 375080
rect 379606 375028 379612 375080
rect 379664 375068 379670 375080
rect 423950 375068 423956 375080
rect 379664 375040 423956 375068
rect 379664 375028 379670 375040
rect 423950 375028 423956 375040
rect 424008 375028 424014 375080
rect 85022 374960 85028 375012
rect 85080 375000 85086 375012
rect 218146 375000 218152 375012
rect 85080 374972 218152 375000
rect 85080 374960 85086 374972
rect 218146 374960 218152 374972
rect 218204 375000 218210 375012
rect 218606 375000 218612 375012
rect 218204 374972 218612 375000
rect 218204 374960 218210 374972
rect 218606 374960 218612 374972
rect 218664 375000 218670 375012
rect 244274 375000 244280 375012
rect 218664 374972 244280 375000
rect 218664 374960 218670 374972
rect 244274 374960 244280 374972
rect 244332 374960 244338 375012
rect 368290 374960 368296 375012
rect 368348 375000 368354 375012
rect 371510 375000 371516 375012
rect 368348 374972 371516 375000
rect 368348 374960 368354 374972
rect 371510 374960 371516 374972
rect 371568 375000 371574 375012
rect 372522 375000 372528 375012
rect 371568 374972 372528 375000
rect 371568 374960 371574 374972
rect 372522 374960 372528 374972
rect 372580 374960 372586 375012
rect 405366 375000 405372 375012
rect 373920 374972 405372 375000
rect 197998 374892 198004 374944
rect 198056 374932 198062 374944
rect 342254 374932 342260 374944
rect 198056 374904 342260 374932
rect 198056 374892 198062 374904
rect 342254 374892 342260 374904
rect 342312 374892 342318 374944
rect 356882 374892 356888 374944
rect 356940 374932 356946 374944
rect 372430 374932 372436 374944
rect 356940 374904 372436 374932
rect 356940 374892 356946 374904
rect 372430 374892 372436 374904
rect 372488 374932 372494 374944
rect 373920 374932 373948 374972
rect 405366 374960 405372 374972
rect 405424 374960 405430 375012
rect 377214 374932 377220 374944
rect 372488 374904 373948 374932
rect 375484 374904 377220 374932
rect 372488 374892 372494 374904
rect 361390 374824 361396 374876
rect 361448 374864 361454 374876
rect 375484 374864 375512 374904
rect 377214 374892 377220 374904
rect 377272 374932 377278 374944
rect 418154 374932 418160 374944
rect 377272 374904 418160 374932
rect 377272 374892 377278 374904
rect 418154 374892 418160 374904
rect 418212 374892 418218 374944
rect 361448 374836 375512 374864
rect 361448 374824 361454 374836
rect 375650 374824 375656 374876
rect 375708 374864 375714 374876
rect 378226 374864 378232 374876
rect 375708 374836 378232 374864
rect 375708 374824 375714 374836
rect 378226 374824 378232 374836
rect 378284 374864 378290 374876
rect 425146 374864 425152 374876
rect 378284 374836 425152 374864
rect 378284 374824 378290 374836
rect 425146 374824 425152 374836
rect 425204 374824 425210 374876
rect 357986 374756 357992 374808
rect 358044 374796 358050 374808
rect 372982 374796 372988 374808
rect 358044 374768 372988 374796
rect 358044 374756 358050 374768
rect 372982 374756 372988 374768
rect 373040 374796 373046 374808
rect 421742 374796 421748 374808
rect 373040 374768 421748 374796
rect 373040 374756 373046 374768
rect 421742 374756 421748 374768
rect 421800 374756 421806 374808
rect 372522 374688 372528 374740
rect 372580 374728 372586 374740
rect 419626 374728 419632 374740
rect 372580 374700 419632 374728
rect 372580 374688 372586 374700
rect 419626 374688 419632 374700
rect 419684 374688 419690 374740
rect 208026 374620 208032 374672
rect 208084 374660 208090 374672
rect 219250 374660 219256 374672
rect 208084 374632 219256 374660
rect 208084 374620 208090 374632
rect 219250 374620 219256 374632
rect 219308 374660 219314 374672
rect 266354 374660 266360 374672
rect 219308 374632 266360 374660
rect 219308 374620 219314 374632
rect 266354 374620 266360 374632
rect 266412 374620 266418 374672
rect 377398 374620 377404 374672
rect 377456 374660 377462 374672
rect 377950 374660 377956 374672
rect 377456 374632 377956 374660
rect 377456 374620 377462 374632
rect 377950 374620 377956 374632
rect 378008 374620 378014 374672
rect 429286 374660 429292 374672
rect 378060 374632 429292 374660
rect 371786 374552 371792 374604
rect 371844 374592 371850 374604
rect 372522 374592 372528 374604
rect 371844 374564 372528 374592
rect 371844 374552 371850 374564
rect 372522 374552 372528 374564
rect 372580 374592 372586 374604
rect 378060 374592 378088 374632
rect 429286 374620 429292 374632
rect 429344 374620 429350 374672
rect 372580 374564 378088 374592
rect 372580 374552 372586 374564
rect 378134 374552 378140 374604
rect 378192 374592 378198 374604
rect 379330 374592 379336 374604
rect 378192 374564 379336 374592
rect 378192 374552 378198 374564
rect 379330 374552 379336 374564
rect 379388 374592 379394 374604
rect 409966 374592 409972 374604
rect 379388 374564 409972 374592
rect 379388 374552 379394 374564
rect 409966 374552 409972 374564
rect 410024 374552 410030 374604
rect 359918 373260 359924 373312
rect 359976 373300 359982 373312
rect 519354 373300 519360 373312
rect 359976 373272 519360 373300
rect 359976 373260 359982 373272
rect 519354 373260 519360 373272
rect 519412 373260 519418 373312
rect 519354 372580 519360 372632
rect 519412 372620 519418 372632
rect 519630 372620 519636 372632
rect 519412 372592 519636 372620
rect 519412 372580 519418 372592
rect 519630 372580 519636 372592
rect 519688 372580 519694 372632
rect 519170 371940 519176 371952
rect 509206 371912 519176 371940
rect 359642 371832 359648 371884
rect 359700 371872 359706 371884
rect 509206 371872 509234 371912
rect 519170 371900 519176 371912
rect 519228 371940 519234 371952
rect 519538 371940 519544 371952
rect 519228 371912 519544 371940
rect 519228 371900 519234 371912
rect 519538 371900 519544 371912
rect 519596 371900 519602 371952
rect 359700 371844 509234 371872
rect 359700 371832 359706 371844
rect 199470 370472 199476 370524
rect 199528 370512 199534 370524
rect 358998 370512 359004 370524
rect 199528 370484 359004 370512
rect 199528 370472 199534 370484
rect 358998 370472 359004 370484
rect 359056 370472 359062 370524
rect 358998 369180 359004 369232
rect 359056 369220 359062 369232
rect 359458 369220 359464 369232
rect 359056 369192 359464 369220
rect 359056 369180 359062 369192
rect 359458 369180 359464 369192
rect 359516 369220 359522 369232
rect 518986 369220 518992 369232
rect 359516 369192 518992 369220
rect 359516 369180 359522 369192
rect 518986 369180 518992 369192
rect 519044 369180 519050 369232
rect 199562 369112 199568 369164
rect 199620 369152 199626 369164
rect 358906 369152 358912 369164
rect 199620 369124 358912 369152
rect 199620 369112 199626 369124
rect 358906 369112 358912 369124
rect 358964 369152 358970 369164
rect 359550 369152 359556 369164
rect 358964 369124 359556 369152
rect 358964 369112 358970 369124
rect 359550 369112 359556 369124
rect 359608 369112 359614 369164
rect 359550 366324 359556 366376
rect 359608 366364 359614 366376
rect 519078 366364 519084 366376
rect 359608 366336 519084 366364
rect 359608 366324 359614 366336
rect 519078 366324 519084 366336
rect 519136 366364 519142 366376
rect 519354 366364 519360 366376
rect 519136 366336 519360 366364
rect 519136 366324 519142 366336
rect 519354 366324 519360 366336
rect 519412 366324 519418 366376
rect 199746 363604 199752 363656
rect 199804 363644 199810 363656
rect 359090 363644 359096 363656
rect 199804 363616 359096 363644
rect 199804 363604 199810 363616
rect 359090 363604 359096 363616
rect 359148 363644 359154 363656
rect 519262 363644 519268 363656
rect 359148 363616 519268 363644
rect 359148 363604 359154 363616
rect 519262 363604 519268 363616
rect 519320 363604 519326 363656
rect 199562 362924 199568 362976
rect 199620 362964 199626 362976
rect 199746 362964 199752 362976
rect 199620 362936 199752 362964
rect 199620 362924 199626 362936
rect 199746 362924 199752 362936
rect 199804 362924 199810 362976
rect 359182 362380 359188 362432
rect 359240 362420 359246 362432
rect 359642 362420 359648 362432
rect 359240 362392 359648 362420
rect 359240 362380 359246 362392
rect 359642 362380 359648 362392
rect 359700 362380 359706 362432
rect 199746 362176 199752 362228
rect 199804 362216 199810 362228
rect 359182 362216 359188 362228
rect 199804 362188 359188 362216
rect 199804 362176 199810 362188
rect 359182 362176 359188 362188
rect 359240 362176 359246 362228
rect 201402 360204 201408 360256
rect 201460 360244 201466 360256
rect 206278 360244 206284 360256
rect 201460 360216 206284 360244
rect 201460 360204 201466 360216
rect 206278 360204 206284 360216
rect 206336 360204 206342 360256
rect 178678 360136 178684 360188
rect 178736 360176 178742 360188
rect 196526 360176 196532 360188
rect 178736 360148 196532 360176
rect 178736 360136 178742 360148
rect 196526 360136 196532 360148
rect 196584 360136 196590 360188
rect 179874 360068 179880 360120
rect 179932 360108 179938 360120
rect 197262 360108 197268 360120
rect 179932 360080 197268 360108
rect 179932 360068 179938 360080
rect 197262 360068 197268 360080
rect 197320 360068 197326 360120
rect 196526 359660 196532 359712
rect 196584 359700 196590 359712
rect 197354 359700 197360 359712
rect 196584 359672 197360 359700
rect 196584 359660 196590 359672
rect 197354 359660 197360 359672
rect 197412 359660 197418 359712
rect 500770 359660 500776 359712
rect 500828 359700 500834 359712
rect 500828 359672 509234 359700
rect 500828 359660 500834 359672
rect 509206 359632 509234 359672
rect 517790 359632 517796 359644
rect 509206 359604 517796 359632
rect 517790 359592 517796 359604
rect 517848 359632 517854 359644
rect 517974 359632 517980 359644
rect 517848 359604 517980 359632
rect 517848 359592 517854 359604
rect 517974 359592 517980 359604
rect 518032 359592 518038 359644
rect 339862 359524 339868 359576
rect 339920 359564 339926 359576
rect 357066 359564 357072 359576
rect 339920 359536 357072 359564
rect 339920 359524 339926 359536
rect 357066 359524 357072 359536
rect 357124 359524 357130 359576
rect 498930 359524 498936 359576
rect 498988 359564 498994 359576
rect 517882 359564 517888 359576
rect 498988 359536 517888 359564
rect 498988 359524 498994 359536
rect 517882 359524 517888 359536
rect 517940 359524 517946 359576
rect 190914 359456 190920 359508
rect 190972 359496 190978 359508
rect 200758 359496 200764 359508
rect 190972 359468 200764 359496
rect 190972 359456 190978 359468
rect 200758 359456 200764 359468
rect 200816 359496 200822 359508
rect 201402 359496 201408 359508
rect 200816 359468 201408 359496
rect 200816 359456 200822 359468
rect 201402 359456 201408 359468
rect 201460 359456 201466 359508
rect 351730 359456 351736 359508
rect 351788 359496 351794 359508
rect 358078 359496 358084 359508
rect 351788 359468 358084 359496
rect 351788 359456 351794 359468
rect 358078 359456 358084 359468
rect 358136 359456 358142 359508
rect 360194 359252 360200 359304
rect 360252 359292 360258 359304
rect 361574 359292 361580 359304
rect 360252 359264 361580 359292
rect 360252 359252 360258 359264
rect 361574 359252 361580 359264
rect 361632 359252 361638 359304
rect 342254 358844 342260 358896
rect 342312 358884 342318 358896
rect 357526 358884 357532 358896
rect 342312 358856 357532 358884
rect 342312 358844 342318 358856
rect 357526 358844 357532 358856
rect 357584 358884 357590 358896
rect 358630 358884 358636 358896
rect 357584 358856 358636 358884
rect 357584 358844 357590 358856
rect 358630 358844 358636 358856
rect 358688 358844 358694 358896
rect 338482 358776 338488 358828
rect 338540 358816 338546 358828
rect 360194 358816 360200 358828
rect 338540 358788 360200 358816
rect 338540 358776 338546 358788
rect 360194 358776 360200 358788
rect 360252 358776 360258 358828
rect 510890 358776 510896 358828
rect 510948 358816 510954 358828
rect 517514 358816 517520 358828
rect 510948 358788 517520 358816
rect 510948 358776 510954 358788
rect 517514 358776 517520 358788
rect 517572 358776 517578 358828
rect 218514 358708 218520 358760
rect 218572 358748 218578 358760
rect 221182 358748 221188 358760
rect 218572 358720 221188 358748
rect 218572 358708 218578 358720
rect 221182 358708 221188 358720
rect 221240 358708 221246 358760
rect 378686 358708 378692 358760
rect 378744 358748 378750 358760
rect 380894 358748 380900 358760
rect 378744 358720 380900 358748
rect 378744 358708 378750 358720
rect 380894 358708 380900 358720
rect 380952 358708 380958 358760
rect 215846 358640 215852 358692
rect 215904 358680 215910 358692
rect 220998 358680 221004 358692
rect 215904 358652 221004 358680
rect 215904 358640 215910 358652
rect 220998 358640 221004 358652
rect 221056 358640 221062 358692
rect 219158 358504 219164 358556
rect 219216 358544 219222 358556
rect 220814 358544 220820 358556
rect 219216 358516 220820 358544
rect 219216 358504 219222 358516
rect 220814 358504 220820 358516
rect 220872 358504 220878 358556
rect 217870 358232 217876 358284
rect 217928 358272 217934 358284
rect 221274 358272 221280 358284
rect 217928 358244 221280 358272
rect 217928 358232 217934 358244
rect 221274 358232 221280 358244
rect 221332 358232 221338 358284
rect 379238 358232 379244 358284
rect 379296 358272 379302 358284
rect 381078 358272 381084 358284
rect 379296 358244 381084 358272
rect 379296 358232 379302 358244
rect 381078 358232 381084 358244
rect 381136 358232 381142 358284
rect 214926 358164 214932 358216
rect 214984 358204 214990 358216
rect 221090 358204 221096 358216
rect 214984 358176 221096 358204
rect 214984 358164 214990 358176
rect 221090 358164 221096 358176
rect 221148 358164 221154 358216
rect 54294 358028 54300 358080
rect 54352 358068 54358 358080
rect 60090 358068 60096 358080
rect 54352 358040 60096 358068
rect 54352 358028 54358 358040
rect 60090 358028 60096 358040
rect 60148 358028 60154 358080
rect 182818 358028 182824 358080
rect 182876 358068 182882 358080
rect 200114 358068 200120 358080
rect 182876 358040 200120 358068
rect 182876 358028 182882 358040
rect 200114 358028 200120 358040
rect 200172 358068 200178 358080
rect 342254 358068 342260 358080
rect 200172 358040 342260 358068
rect 200172 358028 200178 358040
rect 342254 358028 342260 358040
rect 342312 358028 342318 358080
rect 373810 358028 373816 358080
rect 373868 358068 373874 358080
rect 381170 358068 381176 358080
rect 373868 358040 381176 358068
rect 373868 358028 373874 358040
rect 381170 358028 381176 358040
rect 381228 358028 381234 358080
rect 377030 357960 377036 358012
rect 377088 358000 377094 358012
rect 380986 358000 380992 358012
rect 377088 357972 380992 358000
rect 377088 357960 377094 357972
rect 380986 357960 380992 357972
rect 381044 357960 381050 358012
rect 57146 357824 57152 357876
rect 57204 357864 57210 357876
rect 59538 357864 59544 357876
rect 57204 357836 59544 357864
rect 57204 357824 57210 357836
rect 59538 357824 59544 357836
rect 59596 357824 59602 357876
rect 215754 357552 215760 357604
rect 215812 357592 215818 357604
rect 220906 357592 220912 357604
rect 215812 357564 220912 357592
rect 215812 357552 215818 357564
rect 220906 357552 220912 357564
rect 220964 357552 220970 357604
rect 58526 356192 58532 356244
rect 58584 356232 58590 356244
rect 59354 356232 59360 356244
rect 58584 356204 59360 356232
rect 58584 356192 58590 356204
rect 59354 356192 59360 356204
rect 59412 356192 59418 356244
rect 58618 355988 58624 356040
rect 58676 356028 58682 356040
rect 59446 356028 59452 356040
rect 58676 356000 59452 356028
rect 58676 355988 58682 356000
rect 59446 355988 59452 356000
rect 59504 355988 59510 356040
rect 46290 303560 46296 303612
rect 46348 303600 46354 303612
rect 57606 303600 57612 303612
rect 46348 303572 57612 303600
rect 46348 303560 46354 303572
rect 57606 303560 57612 303572
rect 57664 303560 57670 303612
rect 46382 300772 46388 300824
rect 46440 300812 46446 300824
rect 57054 300812 57060 300824
rect 46440 300784 57060 300812
rect 46440 300772 46446 300784
rect 57054 300772 57060 300784
rect 57112 300812 57118 300824
rect 57422 300812 57428 300824
rect 57112 300784 57428 300812
rect 57112 300772 57118 300784
rect 57422 300772 57428 300784
rect 57480 300772 57486 300824
rect 57422 300636 57428 300688
rect 57480 300676 57486 300688
rect 57606 300676 57612 300688
rect 57480 300648 57612 300676
rect 57480 300636 57486 300648
rect 57606 300636 57612 300648
rect 57664 300636 57670 300688
rect 520182 288396 520188 288448
rect 520240 288436 520246 288448
rect 580258 288436 580264 288448
rect 520240 288408 580264 288436
rect 520240 288396 520246 288408
rect 580258 288396 580264 288408
rect 580316 288396 580322 288448
rect 519262 287036 519268 287088
rect 519320 287076 519326 287088
rect 580350 287076 580356 287088
rect 519320 287048 580356 287076
rect 519320 287036 519326 287048
rect 580350 287036 580356 287048
rect 580408 287036 580414 287088
rect 200942 284248 200948 284300
rect 201000 284288 201006 284300
rect 216674 284288 216680 284300
rect 201000 284260 216680 284288
rect 201000 284248 201006 284260
rect 216674 284248 216680 284260
rect 216732 284248 216738 284300
rect 361206 284248 361212 284300
rect 361264 284288 361270 284300
rect 376938 284288 376944 284300
rect 361264 284260 376944 284288
rect 361264 284248 361270 284260
rect 376938 284248 376944 284260
rect 376996 284248 377002 284300
rect 203794 282820 203800 282872
rect 203852 282860 203858 282872
rect 216858 282860 216864 282872
rect 203852 282832 216864 282860
rect 203852 282820 203858 282832
rect 216858 282820 216864 282832
rect 216916 282820 216922 282872
rect 366910 282820 366916 282872
rect 366968 282860 366974 282872
rect 376754 282860 376760 282872
rect 366968 282832 376760 282860
rect 366968 282820 366974 282832
rect 376754 282820 376760 282832
rect 376812 282820 376818 282872
rect 55858 282684 55864 282736
rect 55916 282724 55922 282736
rect 58434 282724 58440 282736
rect 55916 282696 58440 282724
rect 55916 282684 55922 282696
rect 58434 282684 58440 282696
rect 58492 282684 58498 282736
rect 52914 282344 52920 282396
rect 52972 282384 52978 282396
rect 53190 282384 53196 282396
rect 52972 282356 53196 282384
rect 52972 282344 52978 282356
rect 53190 282344 53196 282356
rect 53248 282344 53254 282396
rect 54386 282140 54392 282192
rect 54444 282180 54450 282192
rect 58710 282180 58716 282192
rect 54444 282152 58716 282180
rect 54444 282140 54450 282152
rect 58710 282140 58716 282152
rect 58768 282140 58774 282192
rect 200758 282140 200764 282192
rect 200816 282180 200822 282192
rect 216674 282180 216680 282192
rect 200816 282152 216680 282180
rect 200816 282140 200822 282152
rect 216674 282140 216680 282152
rect 216732 282140 216738 282192
rect 358078 282140 358084 282192
rect 358136 282180 358142 282192
rect 376938 282180 376944 282192
rect 358136 282152 376944 282180
rect 358136 282140 358142 282152
rect 376938 282140 376944 282152
rect 376996 282140 377002 282192
rect 58526 281460 58532 281512
rect 58584 281500 58590 281512
rect 59722 281500 59728 281512
rect 58584 281472 59728 281500
rect 58584 281460 58590 281472
rect 59722 281460 59728 281472
rect 59780 281460 59786 281512
rect 212258 274728 212264 274780
rect 212316 274768 212322 274780
rect 215662 274768 215668 274780
rect 212316 274740 215668 274768
rect 212316 274728 212322 274740
rect 215662 274728 215668 274740
rect 215720 274728 215726 274780
rect 213730 274660 213736 274712
rect 213788 274700 213794 274712
rect 214098 274700 214104 274712
rect 213788 274672 214104 274700
rect 213788 274660 213794 274672
rect 214098 274660 214104 274672
rect 214156 274660 214162 274712
rect 215662 273912 215668 273964
rect 215720 273952 215726 273964
rect 273162 273952 273168 273964
rect 215720 273924 273168 273952
rect 215720 273912 215726 273924
rect 273162 273912 273168 273924
rect 273220 273912 273226 273964
rect 43346 273572 43352 273624
rect 43404 273612 43410 273624
rect 133414 273612 133420 273624
rect 43404 273584 133420 273612
rect 43404 273572 43410 273584
rect 133414 273572 133420 273584
rect 133472 273572 133478 273624
rect 45094 273504 45100 273556
rect 45152 273544 45158 273556
rect 135898 273544 135904 273556
rect 45152 273516 135904 273544
rect 45152 273504 45158 273516
rect 135898 273504 135904 273516
rect 135956 273504 135962 273556
rect 219250 273504 219256 273556
rect 219308 273544 219314 273556
rect 220814 273544 220820 273556
rect 219308 273516 220820 273544
rect 219308 273504 219314 273516
rect 220814 273504 220820 273516
rect 220872 273544 220878 273556
rect 266354 273544 266360 273556
rect 220872 273516 266360 273544
rect 220872 273504 220878 273516
rect 266354 273504 266360 273516
rect 266412 273504 266418 273556
rect 45462 273436 45468 273488
rect 45520 273476 45526 273488
rect 138474 273476 138480 273488
rect 45520 273448 138480 273476
rect 45520 273436 45526 273448
rect 138474 273436 138480 273448
rect 138532 273436 138538 273488
rect 211706 273436 211712 273488
rect 211764 273476 211770 273488
rect 214190 273476 214196 273488
rect 211764 273448 214196 273476
rect 211764 273436 211770 273448
rect 214190 273436 214196 273448
rect 214248 273476 214254 273488
rect 269758 273476 269764 273488
rect 214248 273448 269764 273476
rect 214248 273436 214254 273448
rect 269758 273436 269764 273448
rect 269816 273436 269822 273488
rect 370314 273436 370320 273488
rect 370372 273476 370378 273488
rect 378134 273476 378140 273488
rect 370372 273448 378140 273476
rect 370372 273436 370378 273448
rect 378134 273436 378140 273448
rect 378192 273476 378198 273488
rect 378594 273476 378600 273488
rect 378192 273448 378600 273476
rect 378192 273436 378198 273448
rect 378594 273436 378600 273448
rect 378652 273436 378658 273488
rect 379514 273436 379520 273488
rect 379572 273476 379578 273488
rect 427630 273476 427636 273488
rect 379572 273448 427636 273476
rect 379572 273436 379578 273448
rect 427630 273436 427636 273448
rect 427688 273436 427694 273488
rect 45186 273368 45192 273420
rect 45244 273408 45250 273420
rect 140866 273408 140872 273420
rect 45244 273380 140872 273408
rect 45244 273368 45250 273380
rect 140866 273368 140872 273380
rect 140924 273368 140930 273420
rect 271138 273408 271144 273420
rect 213380 273380 271144 273408
rect 213380 273352 213408 273380
rect 271138 273368 271144 273380
rect 271196 273368 271202 273420
rect 374454 273368 374460 273420
rect 374512 273408 374518 273420
rect 422846 273408 422852 273420
rect 374512 273380 422852 273408
rect 374512 273368 374518 273380
rect 422846 273368 422852 273380
rect 422904 273368 422910 273420
rect 45370 273300 45376 273352
rect 45428 273340 45434 273352
rect 143534 273340 143540 273352
rect 45428 273312 143540 273340
rect 45428 273300 45434 273312
rect 143534 273300 143540 273312
rect 143592 273300 143598 273352
rect 213086 273300 213092 273352
rect 213144 273340 213150 273352
rect 213362 273340 213368 273352
rect 213144 273312 213368 273340
rect 213144 273300 213150 273312
rect 213362 273300 213368 273312
rect 213420 273300 213426 273352
rect 213730 273300 213736 273352
rect 213788 273340 213794 273352
rect 273254 273340 273260 273352
rect 213788 273312 273260 273340
rect 213788 273300 213794 273312
rect 273254 273300 273260 273312
rect 273312 273300 273318 273352
rect 366726 273300 366732 273352
rect 366784 273340 366790 273352
rect 421098 273340 421104 273352
rect 366784 273312 421104 273340
rect 366784 273300 366790 273312
rect 421098 273300 421104 273312
rect 421156 273300 421162 273352
rect 45278 273232 45284 273284
rect 45336 273272 45342 273284
rect 145926 273272 145932 273284
rect 45336 273244 145932 273272
rect 45336 273232 45342 273244
rect 145926 273232 145932 273244
rect 145984 273232 145990 273284
rect 206738 273232 206744 273284
rect 206796 273272 206802 273284
rect 283466 273272 283472 273284
rect 206796 273244 283472 273272
rect 206796 273232 206802 273244
rect 283466 273232 283472 273244
rect 283524 273232 283530 273284
rect 370866 273232 370872 273284
rect 370924 273272 370930 273284
rect 445938 273272 445944 273284
rect 370924 273244 445944 273272
rect 370924 273232 370930 273244
rect 445938 273232 445944 273244
rect 445996 273232 446002 273284
rect 42334 273164 42340 273216
rect 42392 273204 42398 273216
rect 46014 273204 46020 273216
rect 42392 273176 46020 273204
rect 42392 273164 42398 273176
rect 46014 273164 46020 273176
rect 46072 273164 46078 273216
rect 378594 273164 378600 273216
rect 378652 273204 378658 273216
rect 425238 273204 425244 273216
rect 378652 273176 425244 273204
rect 378652 273164 378658 273176
rect 425238 273164 425244 273176
rect 425296 273164 425302 273216
rect 212350 273096 212356 273148
rect 212408 273136 212414 273148
rect 285950 273136 285956 273148
rect 212408 273108 285956 273136
rect 212408 273096 212414 273108
rect 285950 273096 285956 273108
rect 286008 273096 286014 273148
rect 369578 273096 369584 273148
rect 369636 273136 369642 273148
rect 423398 273136 423404 273148
rect 369636 273108 423404 273136
rect 369636 273096 369642 273108
rect 423398 273096 423404 273108
rect 423456 273096 423462 273148
rect 209314 273028 209320 273080
rect 209372 273068 209378 273080
rect 288158 273068 288164 273080
rect 209372 273040 288164 273068
rect 209372 273028 209378 273040
rect 288158 273028 288164 273040
rect 288216 273028 288222 273080
rect 356790 273028 356796 273080
rect 356848 273068 356854 273080
rect 425974 273068 425980 273080
rect 356848 273040 425980 273068
rect 356848 273028 356854 273040
rect 425974 273028 425980 273040
rect 426032 273028 426038 273080
rect 216306 272960 216312 273012
rect 216364 273000 216370 273012
rect 298462 273000 298468 273012
rect 216364 272972 298468 273000
rect 216364 272960 216370 272972
rect 298462 272960 298468 272972
rect 298520 272960 298526 273012
rect 358446 272960 358452 273012
rect 358504 273000 358510 273012
rect 428182 273000 428188 273012
rect 358504 272972 428188 273000
rect 358504 272960 358510 272972
rect 428182 272960 428188 272972
rect 428240 272960 428246 273012
rect 210878 272892 210884 272944
rect 210936 272932 210942 272944
rect 295886 272932 295892 272944
rect 210936 272904 295892 272932
rect 210936 272892 210942 272904
rect 295886 272892 295892 272904
rect 295944 272892 295950 272944
rect 372338 272892 372344 272944
rect 372396 272932 372402 272944
rect 468478 272932 468484 272944
rect 372396 272904 468484 272932
rect 372396 272892 372402 272904
rect 468478 272892 468484 272904
rect 468536 272892 468542 272944
rect 42426 272824 42432 272876
rect 42484 272864 42490 272876
rect 60826 272864 60832 272876
rect 42484 272836 60832 272864
rect 42484 272824 42490 272836
rect 60826 272824 60832 272836
rect 60884 272824 60890 272876
rect 202414 272824 202420 272876
rect 202472 272864 202478 272876
rect 290918 272864 290924 272876
rect 202472 272836 290924 272864
rect 202472 272824 202478 272836
rect 290918 272824 290924 272836
rect 290976 272824 290982 272876
rect 373442 272824 373448 272876
rect 373500 272864 373506 272876
rect 478414 272864 478420 272876
rect 373500 272836 478420 272864
rect 373500 272824 373506 272836
rect 478414 272824 478420 272836
rect 478472 272824 478478 272876
rect 48130 272756 48136 272808
rect 48188 272796 48194 272808
rect 77110 272796 77116 272808
rect 48188 272768 77116 272796
rect 48188 272756 48194 272768
rect 77110 272756 77116 272768
rect 77168 272756 77174 272808
rect 203702 272756 203708 272808
rect 203760 272796 203766 272808
rect 293310 272796 293316 272808
rect 203760 272768 293316 272796
rect 203760 272756 203766 272768
rect 293310 272756 293316 272768
rect 293368 272756 293374 272808
rect 363966 272756 363972 272808
rect 364024 272796 364030 272808
rect 470870 272796 470876 272808
rect 364024 272768 470876 272796
rect 364024 272756 364030 272768
rect 470870 272756 470876 272768
rect 470928 272756 470934 272808
rect 50430 272688 50436 272740
rect 50488 272728 50494 272740
rect 90726 272728 90732 272740
rect 50488 272700 90732 272728
rect 50488 272688 50494 272700
rect 90726 272688 90732 272700
rect 90784 272688 90790 272740
rect 207842 272688 207848 272740
rect 207900 272728 207906 272740
rect 300854 272728 300860 272740
rect 207900 272700 300860 272728
rect 207900 272688 207906 272700
rect 300854 272688 300860 272700
rect 300912 272688 300918 272740
rect 365346 272688 365352 272740
rect 365404 272728 365410 272740
rect 473446 272728 473452 272740
rect 365404 272700 473452 272728
rect 365404 272688 365410 272700
rect 473446 272688 473452 272700
rect 473504 272688 473510 272740
rect 48958 272620 48964 272672
rect 49016 272660 49022 272672
rect 50246 272660 50252 272672
rect 49016 272632 50252 272660
rect 49016 272620 49022 272632
rect 50246 272620 50252 272632
rect 50304 272620 50310 272672
rect 51626 272620 51632 272672
rect 51684 272660 51690 272672
rect 93670 272660 93676 272672
rect 51684 272632 93676 272660
rect 51684 272620 51690 272632
rect 93670 272620 93676 272632
rect 93728 272620 93734 272672
rect 205266 272620 205272 272672
rect 205324 272660 205330 272672
rect 303430 272660 303436 272672
rect 205324 272632 303436 272660
rect 205324 272620 205330 272632
rect 303430 272620 303436 272632
rect 303488 272620 303494 272672
rect 368198 272620 368204 272672
rect 368256 272660 368262 272672
rect 480806 272660 480812 272672
rect 368256 272632 480812 272660
rect 368256 272620 368262 272632
rect 480806 272620 480812 272632
rect 480864 272620 480870 272672
rect 48038 272552 48044 272604
rect 48096 272592 48102 272604
rect 95878 272592 95884 272604
rect 48096 272564 95884 272592
rect 48096 272552 48102 272564
rect 95878 272552 95884 272564
rect 95936 272552 95942 272604
rect 206554 272552 206560 272604
rect 206612 272592 206618 272604
rect 310974 272592 310980 272604
rect 206612 272564 310980 272592
rect 206612 272552 206618 272564
rect 310974 272552 310980 272564
rect 311032 272552 311038 272604
rect 362586 272552 362592 272604
rect 362644 272592 362650 272604
rect 475838 272592 475844 272604
rect 362644 272564 475844 272592
rect 362644 272552 362650 272564
rect 475838 272552 475844 272564
rect 475896 272552 475902 272604
rect 50522 272484 50528 272536
rect 50580 272524 50586 272536
rect 98454 272524 98460 272536
rect 50580 272496 98460 272524
rect 50580 272484 50586 272496
rect 98454 272484 98460 272496
rect 98512 272484 98518 272536
rect 107470 272484 107476 272536
rect 107528 272524 107534 272536
rect 196894 272524 196900 272536
rect 107528 272496 196900 272524
rect 107528 272484 107534 272496
rect 196894 272484 196900 272496
rect 196952 272484 196958 272536
rect 200850 272484 200856 272536
rect 200908 272524 200914 272536
rect 320910 272524 320916 272536
rect 200908 272496 320916 272524
rect 200908 272484 200914 272496
rect 320910 272484 320916 272496
rect 320968 272484 320974 272536
rect 361114 272484 361120 272536
rect 361172 272524 361178 272536
rect 485958 272524 485964 272536
rect 361172 272496 485964 272524
rect 361172 272484 361178 272496
rect 485958 272484 485964 272496
rect 486016 272484 486022 272536
rect 49050 272416 49056 272468
rect 49108 272456 49114 272468
rect 50062 272456 50068 272468
rect 49108 272428 50068 272456
rect 49108 272416 49114 272428
rect 50062 272416 50068 272428
rect 50120 272416 50126 272468
rect 76006 272456 76012 272468
rect 55186 272428 76012 272456
rect 46658 272348 46664 272400
rect 46716 272388 46722 272400
rect 55186 272388 55214 272428
rect 76006 272416 76012 272428
rect 76064 272416 76070 272468
rect 46716 272360 55214 272388
rect 46716 272348 46722 272360
rect 58618 272348 58624 272400
rect 58676 272388 58682 272400
rect 59446 272388 59452 272400
rect 58676 272360 59452 272388
rect 58676 272348 58682 272360
rect 59446 272348 59452 272360
rect 59504 272348 59510 272400
rect 62114 272348 62120 272400
rect 62172 272388 62178 272400
rect 94406 272388 94412 272400
rect 62172 272360 94412 272388
rect 62172 272348 62178 272360
rect 94406 272348 94412 272360
rect 94464 272348 94470 272400
rect 50062 272280 50068 272332
rect 50120 272320 50126 272332
rect 82998 272320 83004 272332
rect 50120 272292 83004 272320
rect 50120 272280 50126 272292
rect 82998 272280 83004 272292
rect 83056 272280 83062 272332
rect 374362 272280 374368 272332
rect 374420 272320 374426 272332
rect 375098 272320 375104 272332
rect 374420 272292 375104 272320
rect 374420 272280 374426 272292
rect 375098 272280 375104 272292
rect 375156 272280 375162 272332
rect 58434 272212 58440 272264
rect 58492 272252 58498 272264
rect 60734 272252 60740 272264
rect 58492 272224 60740 272252
rect 58492 272212 58498 272224
rect 60734 272212 60740 272224
rect 60792 272252 60798 272264
rect 100754 272252 100760 272264
rect 60792 272224 100760 272252
rect 60792 272212 60798 272224
rect 100754 272212 100760 272224
rect 100812 272212 100818 272264
rect 46474 272144 46480 272196
rect 46532 272184 46538 272196
rect 51442 272184 51448 272196
rect 46532 272156 51448 272184
rect 46532 272144 46538 272156
rect 51442 272144 51448 272156
rect 51500 272184 51506 272196
rect 51500 272156 55214 272184
rect 51500 272144 51506 272156
rect 46566 272076 46572 272128
rect 46624 272116 46630 272128
rect 48958 272116 48964 272128
rect 46624 272088 48964 272116
rect 46624 272076 46630 272088
rect 48958 272076 48964 272088
rect 49016 272076 49022 272128
rect 55186 272116 55214 272156
rect 58710 272144 58716 272196
rect 58768 272184 58774 272196
rect 60918 272184 60924 272196
rect 58768 272156 60924 272184
rect 58768 272144 58774 272156
rect 60918 272144 60924 272156
rect 60976 272184 60982 272196
rect 102134 272184 102140 272196
rect 60976 272156 102140 272184
rect 60976 272144 60982 272156
rect 102134 272144 102140 272156
rect 102192 272144 102198 272196
rect 95970 272116 95976 272128
rect 55186 272088 95976 272116
rect 95970 272076 95976 272088
rect 96028 272076 96034 272128
rect 371786 272076 371792 272128
rect 371844 272116 371850 272128
rect 373074 272116 373080 272128
rect 371844 272088 373080 272116
rect 371844 272076 371850 272088
rect 373074 272076 373080 272088
rect 373132 272116 373138 272128
rect 433334 272116 433340 272128
rect 373132 272088 433340 272116
rect 373132 272076 373138 272088
rect 433334 272076 433340 272088
rect 433392 272076 433398 272128
rect 52730 272008 52736 272060
rect 52788 272048 52794 272060
rect 53282 272048 53288 272060
rect 52788 272020 53288 272048
rect 52788 272008 52794 272020
rect 53282 272008 53288 272020
rect 53340 272008 53346 272060
rect 60826 272008 60832 272060
rect 60884 272048 60890 272060
rect 104894 272048 104900 272060
rect 60884 272020 104900 272048
rect 60884 272008 60890 272020
rect 104894 272008 104900 272020
rect 104952 272008 104958 272060
rect 373902 272008 373908 272060
rect 373960 272048 373966 272060
rect 379606 272048 379612 272060
rect 373960 272020 379612 272048
rect 373960 272008 373966 272020
rect 379606 272008 379612 272020
rect 379664 272008 379670 272060
rect 396718 272008 396724 272060
rect 396776 272048 396782 272060
rect 415854 272048 415860 272060
rect 396776 272020 415860 272048
rect 396776 272008 396782 272020
rect 415854 272008 415860 272020
rect 415912 272008 415918 272060
rect 48958 271940 48964 271992
rect 49016 271980 49022 271992
rect 97994 271980 98000 271992
rect 49016 271952 98000 271980
rect 49016 271940 49022 271952
rect 97994 271940 98000 271952
rect 98052 271940 98058 271992
rect 370406 271940 370412 271992
rect 370464 271980 370470 271992
rect 372338 271980 372344 271992
rect 370464 271952 372344 271980
rect 370464 271940 370470 271952
rect 372338 271940 372344 271952
rect 372396 271980 372402 271992
rect 430574 271980 430580 271992
rect 372396 271952 430580 271980
rect 372396 271940 372402 271952
rect 430574 271940 430580 271952
rect 430632 271940 430638 271992
rect 48222 271872 48228 271924
rect 48280 271912 48286 271924
rect 107470 271912 107476 271924
rect 48280 271884 107476 271912
rect 48280 271872 48286 271884
rect 107470 271872 107476 271884
rect 107528 271872 107534 271924
rect 114462 271872 114468 271924
rect 114520 271912 114526 271924
rect 127618 271912 127624 271924
rect 114520 271884 127624 271912
rect 114520 271872 114526 271884
rect 127618 271872 127624 271884
rect 127676 271872 127682 271924
rect 215846 271872 215852 271924
rect 215904 271912 215910 271924
rect 216306 271912 216312 271924
rect 215904 271884 216312 271912
rect 215904 271872 215910 271884
rect 216306 271872 216312 271884
rect 216364 271912 216370 271924
rect 276014 271912 276020 271924
rect 216364 271884 276020 271912
rect 216364 271872 216370 271884
rect 276014 271872 276020 271884
rect 276072 271872 276078 271924
rect 356790 271872 356796 271924
rect 356848 271912 356854 271924
rect 359366 271912 359372 271924
rect 356848 271884 359372 271912
rect 356848 271872 356854 271884
rect 359366 271872 359372 271884
rect 359424 271872 359430 271924
rect 360286 271912 360292 271924
rect 359476 271884 360292 271912
rect 43438 271804 43444 271856
rect 43496 271844 43502 271856
rect 129734 271844 129740 271856
rect 43496 271816 129740 271844
rect 43496 271804 43502 271816
rect 129734 271804 129740 271816
rect 129792 271804 129798 271856
rect 154482 271804 154488 271856
rect 154540 271844 154546 271856
rect 201678 271844 201684 271856
rect 154540 271816 201684 271844
rect 154540 271804 154546 271816
rect 201678 271804 201684 271816
rect 201736 271804 201742 271856
rect 343542 271804 343548 271856
rect 343600 271844 343606 271856
rect 358630 271844 358636 271856
rect 343600 271816 358636 271844
rect 343600 271804 343606 271816
rect 358630 271804 358636 271816
rect 358688 271844 358694 271856
rect 359476 271844 359504 271884
rect 360286 271872 360292 271884
rect 360344 271872 360350 271924
rect 425698 271872 425704 271924
rect 425756 271912 425762 271924
rect 427814 271912 427820 271924
rect 425756 271884 427820 271912
rect 425756 271872 425762 271884
rect 427814 271872 427820 271884
rect 427872 271872 427878 271924
rect 358688 271816 359504 271844
rect 358688 271804 358694 271816
rect 369486 271804 369492 271856
rect 369544 271844 369550 271856
rect 458174 271844 458180 271856
rect 369544 271816 458180 271844
rect 369544 271804 369550 271816
rect 458174 271804 458180 271816
rect 458232 271804 458238 271856
rect 517698 271804 517704 271856
rect 517756 271844 517762 271856
rect 517882 271844 517888 271856
rect 517756 271816 517888 271844
rect 517756 271804 517762 271816
rect 517882 271804 517888 271816
rect 517940 271804 517946 271856
rect 42242 271736 42248 271788
rect 42300 271776 42306 271788
rect 123202 271776 123208 271788
rect 42300 271748 123208 271776
rect 42300 271736 42306 271748
rect 123202 271736 123208 271748
rect 123260 271736 123266 271788
rect 158622 271736 158628 271788
rect 158680 271776 158686 271788
rect 205634 271776 205640 271788
rect 158680 271748 205640 271776
rect 158680 271736 158686 271748
rect 205634 271736 205640 271748
rect 205692 271736 205698 271788
rect 212166 271736 212172 271788
rect 212224 271776 212230 271788
rect 307754 271776 307760 271788
rect 212224 271748 307760 271776
rect 212224 271736 212230 271748
rect 307754 271736 307760 271748
rect 307812 271736 307818 271788
rect 368014 271736 368020 271788
rect 368072 271776 368078 271788
rect 455782 271776 455788 271788
rect 368072 271748 455788 271776
rect 368072 271736 368078 271748
rect 455782 271736 455788 271748
rect 455840 271736 455846 271788
rect 42518 271668 42524 271720
rect 42576 271708 42582 271720
rect 52454 271708 52460 271720
rect 42576 271680 52460 271708
rect 42576 271668 42582 271680
rect 52454 271668 52460 271680
rect 52512 271708 52518 271720
rect 52822 271708 52828 271720
rect 52512 271680 52828 271708
rect 52512 271668 52518 271680
rect 52822 271668 52828 271680
rect 52880 271668 52886 271720
rect 54294 271668 54300 271720
rect 54352 271708 54358 271720
rect 125594 271708 125600 271720
rect 54352 271680 125600 271708
rect 54352 271668 54358 271680
rect 125594 271668 125600 271680
rect 125652 271668 125658 271720
rect 151354 271668 151360 271720
rect 151412 271708 151418 271720
rect 197630 271708 197636 271720
rect 151412 271680 197636 271708
rect 151412 271668 151418 271680
rect 197630 271668 197636 271680
rect 197688 271668 197694 271720
rect 202138 271668 202144 271720
rect 202196 271708 202202 271720
rect 270494 271708 270500 271720
rect 202196 271680 270500 271708
rect 202196 271668 202202 271680
rect 270494 271668 270500 271680
rect 270552 271668 270558 271720
rect 363874 271668 363880 271720
rect 363932 271708 363938 271720
rect 449894 271708 449900 271720
rect 363932 271680 449900 271708
rect 363932 271668 363938 271680
rect 449894 271668 449900 271680
rect 449952 271668 449958 271720
rect 57146 271600 57152 271652
rect 57204 271640 57210 271652
rect 128354 271640 128360 271652
rect 57204 271612 128360 271640
rect 57204 271600 57210 271612
rect 128354 271600 128360 271612
rect 128412 271600 128418 271652
rect 157242 271600 157248 271652
rect 157300 271640 157306 271652
rect 202874 271640 202880 271652
rect 157300 271612 202880 271640
rect 157300 271600 157306 271612
rect 202874 271600 202880 271612
rect 202932 271600 202938 271652
rect 214742 271600 214748 271652
rect 214800 271640 214806 271652
rect 280154 271640 280160 271652
rect 214800 271612 280160 271640
rect 214800 271600 214806 271612
rect 280154 271600 280160 271612
rect 280212 271600 280218 271652
rect 370774 271600 370780 271652
rect 370832 271640 370838 271652
rect 452654 271640 452660 271652
rect 370832 271612 452660 271640
rect 370832 271600 370838 271612
rect 452654 271600 452660 271612
rect 452712 271600 452718 271652
rect 54662 271532 54668 271584
rect 54720 271572 54726 271584
rect 120074 271572 120080 271584
rect 54720 271544 120080 271572
rect 54720 271532 54726 271544
rect 120074 271532 120080 271544
rect 120132 271532 120138 271584
rect 161290 271532 161296 271584
rect 161348 271572 161354 271584
rect 204254 271572 204260 271584
rect 161348 271544 204260 271572
rect 161348 271532 161354 271544
rect 204254 271532 204260 271544
rect 204312 271532 204318 271584
rect 216214 271532 216220 271584
rect 216272 271572 216278 271584
rect 276014 271572 276020 271584
rect 216272 271544 276020 271572
rect 216272 271532 216278 271544
rect 276014 271532 276020 271544
rect 276072 271532 276078 271584
rect 368106 271532 368112 271584
rect 368164 271572 368170 271584
rect 442994 271572 443000 271584
rect 368164 271544 443000 271572
rect 368164 271532 368170 271544
rect 442994 271532 443000 271544
rect 443052 271532 443058 271584
rect 53098 271464 53104 271516
rect 53156 271504 53162 271516
rect 115934 271504 115940 271516
rect 53156 271476 115940 271504
rect 53156 271464 53162 271476
rect 115934 271464 115940 271476
rect 115992 271464 115998 271516
rect 164142 271464 164148 271516
rect 164200 271504 164206 271516
rect 197722 271504 197728 271516
rect 164200 271476 197728 271504
rect 164200 271464 164206 271476
rect 197722 271464 197728 271476
rect 197780 271464 197786 271516
rect 205174 271464 205180 271516
rect 205232 271504 205238 271516
rect 263594 271504 263600 271516
rect 205232 271476 263600 271504
rect 205232 271464 205238 271476
rect 263594 271464 263600 271476
rect 263652 271464 263658 271516
rect 372246 271464 372252 271516
rect 372304 271504 372310 271516
rect 447134 271504 447140 271516
rect 372304 271476 447140 271504
rect 372304 271464 372310 271476
rect 447134 271464 447140 271476
rect 447192 271464 447198 271516
rect 46750 271396 46756 271448
rect 46808 271436 46814 271448
rect 53834 271436 53840 271448
rect 46808 271408 53840 271436
rect 46808 271396 46814 271408
rect 53834 271396 53840 271408
rect 53892 271396 53898 271448
rect 54754 271396 54760 271448
rect 54812 271436 54818 271448
rect 117314 271436 117320 271448
rect 54812 271408 117320 271436
rect 54812 271396 54818 271408
rect 117314 271396 117320 271408
rect 117372 271396 117378 271448
rect 166902 271396 166908 271448
rect 166960 271436 166966 271448
rect 166960 271408 180794 271436
rect 166960 271396 166966 271408
rect 53190 271328 53196 271380
rect 53248 271368 53254 271380
rect 113174 271368 113180 271380
rect 53248 271340 113180 271368
rect 53248 271328 53254 271340
rect 113174 271328 113180 271340
rect 113232 271328 113238 271380
rect 180766 271368 180794 271408
rect 196618 271396 196624 271448
rect 196676 271436 196682 271448
rect 197814 271436 197820 271448
rect 196676 271408 197820 271436
rect 196676 271396 196682 271408
rect 197814 271396 197820 271408
rect 197872 271396 197878 271448
rect 219066 271396 219072 271448
rect 219124 271436 219130 271448
rect 277946 271436 277952 271448
rect 219124 271408 277952 271436
rect 219124 271396 219130 271408
rect 277946 271396 277952 271408
rect 278004 271396 278010 271448
rect 361022 271396 361028 271448
rect 361080 271436 361086 271448
rect 426986 271436 426992 271448
rect 361080 271408 426992 271436
rect 361080 271396 361086 271408
rect 426986 271396 426992 271408
rect 427044 271396 427050 271448
rect 427078 271396 427084 271448
rect 427136 271436 427142 271448
rect 432046 271436 432052 271448
rect 427136 271408 432052 271436
rect 427136 271396 427142 271408
rect 432046 271396 432052 271408
rect 432104 271396 432110 271448
rect 200298 271368 200304 271380
rect 180766 271340 200304 271368
rect 200298 271328 200304 271340
rect 200356 271328 200362 271380
rect 203610 271328 203616 271380
rect 203668 271368 203674 271380
rect 260834 271368 260840 271380
rect 203668 271340 260840 271368
rect 203668 271328 203674 271340
rect 260834 271328 260840 271340
rect 260892 271328 260898 271380
rect 362494 271328 362500 271380
rect 362552 271368 362558 271380
rect 434714 271368 434720 271380
rect 362552 271340 434720 271368
rect 362552 271328 362558 271340
rect 434714 271328 434720 271340
rect 434772 271328 434778 271380
rect 503622 271328 503628 271380
rect 503680 271368 503686 271380
rect 517606 271368 517612 271380
rect 503680 271340 517612 271368
rect 503680 271328 503686 271340
rect 517606 271328 517612 271340
rect 517664 271328 517670 271380
rect 51534 271260 51540 271312
rect 51592 271300 51598 271312
rect 110414 271300 110420 271312
rect 51592 271272 110420 271300
rect 51592 271260 51598 271272
rect 110414 271260 110420 271272
rect 110472 271260 110478 271312
rect 197906 271260 197912 271312
rect 197964 271300 197970 271312
rect 200114 271300 200120 271312
rect 197964 271272 200120 271300
rect 197964 271260 197970 271272
rect 200114 271260 200120 271272
rect 200172 271260 200178 271312
rect 210694 271260 210700 271312
rect 210752 271300 210758 271312
rect 267826 271300 267832 271312
rect 210752 271272 267832 271300
rect 210752 271260 210758 271272
rect 267826 271260 267832 271272
rect 267884 271260 267890 271312
rect 343542 271260 343548 271312
rect 343600 271300 343606 271312
rect 356790 271300 356796 271312
rect 343600 271272 356796 271300
rect 343600 271260 343606 271272
rect 356790 271260 356796 271272
rect 356848 271260 356854 271312
rect 366818 271260 366824 271312
rect 366876 271300 366882 271312
rect 437474 271300 437480 271312
rect 366876 271272 437480 271300
rect 366876 271260 366882 271272
rect 437474 271260 437480 271272
rect 437532 271260 437538 271312
rect 52914 271192 52920 271244
rect 52972 271232 52978 271244
rect 107654 271232 107660 271244
rect 52972 271204 107660 271232
rect 52972 271192 52978 271204
rect 107654 271192 107660 271204
rect 107712 271192 107718 271244
rect 183462 271192 183468 271244
rect 183520 271232 183526 271244
rect 197446 271232 197452 271244
rect 183520 271204 197452 271232
rect 183520 271192 183526 271204
rect 197446 271192 197452 271204
rect 197504 271232 197510 271244
rect 197998 271232 198004 271244
rect 197504 271204 198004 271232
rect 197504 271192 197510 271204
rect 197998 271192 198004 271204
rect 198056 271192 198062 271244
rect 209406 271192 209412 271244
rect 209464 271232 209470 271244
rect 264974 271232 264980 271244
rect 209464 271204 264980 271232
rect 209464 271192 209470 271204
rect 264974 271192 264980 271204
rect 265032 271192 265038 271244
rect 278682 271192 278688 271244
rect 278740 271232 278746 271244
rect 357434 271232 357440 271244
rect 278740 271204 357440 271232
rect 278740 271192 278746 271204
rect 357434 271192 357440 271204
rect 357492 271192 357498 271244
rect 373626 271192 373632 271244
rect 373684 271232 373690 271244
rect 440234 271232 440240 271244
rect 373684 271204 440240 271232
rect 373684 271192 373690 271204
rect 440234 271192 440240 271204
rect 440292 271192 440298 271244
rect 503622 271192 503628 271244
rect 503680 271232 503686 271244
rect 517882 271232 517888 271244
rect 503680 271204 517888 271232
rect 503680 271192 503686 271204
rect 517882 271192 517888 271204
rect 517940 271192 517946 271244
rect 51810 271124 51816 271176
rect 51868 271164 51874 271176
rect 104894 271164 104900 271176
rect 51868 271136 104900 271164
rect 51868 271124 51874 271136
rect 104894 271124 104900 271136
rect 104952 271124 104958 271176
rect 127618 271124 127624 271176
rect 127676 271164 127682 271176
rect 196618 271164 196624 271176
rect 127676 271136 196624 271164
rect 127676 271124 127682 271136
rect 196618 271124 196624 271136
rect 196676 271124 196682 271176
rect 206646 271124 206652 271176
rect 206704 271164 206710 271176
rect 258258 271164 258264 271176
rect 206704 271136 258264 271164
rect 206704 271124 206710 271136
rect 258258 271124 258264 271136
rect 258316 271124 258322 271176
rect 275922 271124 275928 271176
rect 275980 271164 275986 271176
rect 356606 271164 356612 271176
rect 275980 271136 356612 271164
rect 275980 271124 275986 271136
rect 356606 271124 356612 271136
rect 356664 271164 356670 271176
rect 356790 271164 356796 271176
rect 356664 271136 356796 271164
rect 356664 271124 356670 271136
rect 356790 271124 356796 271136
rect 356848 271124 356854 271176
rect 358538 271124 358544 271176
rect 358596 271164 358602 271176
rect 416038 271164 416044 271176
rect 358596 271136 416044 271164
rect 358596 271124 358602 271136
rect 416038 271124 416044 271136
rect 416096 271124 416102 271176
rect 426986 271124 426992 271176
rect 427044 271164 427050 271176
rect 433334 271164 433340 271176
rect 427044 271136 433340 271164
rect 427044 271124 427050 271136
rect 433334 271124 433340 271136
rect 433392 271124 433398 271176
rect 440142 271124 440148 271176
rect 440200 271164 440206 271176
rect 516594 271164 516600 271176
rect 440200 271136 516600 271164
rect 440200 271124 440206 271136
rect 516594 271124 516600 271136
rect 516652 271124 516658 271176
rect 51902 271056 51908 271108
rect 51960 271096 51966 271108
rect 103514 271096 103520 271108
rect 51960 271068 103520 271096
rect 51960 271056 51966 271068
rect 103514 271056 103520 271068
rect 103572 271056 103578 271108
rect 209222 271056 209228 271108
rect 209280 271096 209286 271108
rect 255314 271096 255320 271108
rect 209280 271068 255320 271096
rect 209280 271056 209286 271068
rect 255314 271056 255320 271068
rect 255372 271056 255378 271108
rect 379146 271056 379152 271108
rect 379204 271096 379210 271108
rect 418154 271096 418160 271108
rect 379204 271068 418160 271096
rect 379204 271056 379210 271068
rect 418154 271056 418160 271068
rect 418212 271056 418218 271108
rect 50338 270988 50344 271040
rect 50396 271028 50402 271040
rect 100754 271028 100760 271040
rect 50396 271000 100760 271028
rect 50396 270988 50402 271000
rect 100754 270988 100760 271000
rect 100812 270988 100818 271040
rect 210786 270988 210792 271040
rect 210844 271028 210850 271040
rect 252554 271028 252560 271040
rect 210844 271000 252560 271028
rect 210844 270988 210850 271000
rect 252554 270988 252560 271000
rect 252612 270988 252618 271040
rect 374914 270988 374920 271040
rect 374972 271028 374978 271040
rect 412726 271028 412732 271040
rect 374972 271000 412732 271028
rect 374972 270988 374978 271000
rect 412726 270988 412732 271000
rect 412784 270988 412790 271040
rect 54570 270920 54576 270972
rect 54628 270960 54634 270972
rect 88334 270960 88340 270972
rect 54628 270932 88340 270960
rect 54628 270920 54634 270932
rect 88334 270920 88340 270932
rect 88392 270920 88398 270972
rect 214834 270920 214840 270972
rect 214892 270960 214898 270972
rect 247034 270960 247040 270972
rect 214892 270932 247040 270960
rect 214892 270920 214898 270932
rect 247034 270920 247040 270932
rect 247092 270920 247098 270972
rect 374822 270920 374828 270972
rect 374880 270960 374886 270972
rect 409874 270960 409880 270972
rect 374880 270932 409880 270960
rect 374880 270920 374886 270932
rect 409874 270920 409880 270932
rect 409932 270920 409938 270972
rect 213270 270852 213276 270904
rect 213328 270892 213334 270904
rect 313274 270892 313280 270904
rect 213328 270864 313280 270892
rect 213328 270852 213334 270864
rect 313274 270852 313280 270864
rect 313332 270852 313338 270904
rect 183462 270512 183468 270564
rect 183520 270552 183526 270564
rect 197722 270552 197728 270564
rect 183520 270524 197728 270552
rect 183520 270512 183526 270524
rect 197722 270512 197728 270524
rect 197780 270552 197786 270564
rect 197906 270552 197912 270564
rect 197780 270524 197912 270552
rect 197780 270512 197786 270524
rect 197906 270512 197912 270524
rect 197964 270512 197970 270564
rect 47946 270444 47952 270496
rect 48004 270484 48010 270496
rect 147674 270484 147680 270496
rect 48004 270456 147680 270484
rect 48004 270444 48010 270456
rect 147674 270444 147680 270456
rect 147732 270444 147738 270496
rect 212994 270444 213000 270496
rect 213052 270484 213058 270496
rect 213454 270484 213460 270496
rect 213052 270456 213460 270484
rect 213052 270444 213058 270456
rect 213454 270444 213460 270456
rect 213512 270444 213518 270496
rect 219802 270484 219808 270496
rect 219406 270456 219808 270484
rect 53190 270376 53196 270428
rect 53248 270416 53254 270428
rect 86954 270416 86960 270428
rect 53248 270388 86960 270416
rect 53248 270376 53254 270388
rect 86954 270376 86960 270388
rect 87012 270376 87018 270428
rect 216858 270376 216864 270428
rect 216916 270416 216922 270428
rect 219406 270416 219434 270456
rect 219802 270444 219808 270456
rect 219860 270484 219866 270496
rect 247034 270484 247040 270496
rect 219860 270456 247040 270484
rect 219860 270444 219866 270456
rect 247034 270444 247040 270456
rect 247092 270444 247098 270496
rect 280062 270444 280068 270496
rect 280120 270484 280126 270496
rect 356606 270484 356612 270496
rect 280120 270456 356612 270484
rect 280120 270444 280126 270456
rect 356606 270444 356612 270456
rect 356664 270484 356670 270496
rect 357158 270484 357164 270496
rect 356664 270456 357164 270484
rect 356664 270444 356670 270456
rect 357158 270444 357164 270456
rect 357216 270444 357222 270496
rect 365530 270444 365536 270496
rect 365588 270484 365594 270496
rect 368290 270484 368296 270496
rect 365588 270456 368296 270484
rect 365588 270444 365594 270456
rect 368290 270444 368296 270456
rect 368348 270444 368354 270496
rect 377214 270444 377220 270496
rect 377272 270484 377278 270496
rect 377490 270484 377496 270496
rect 377272 270456 377496 270484
rect 377272 270444 377278 270456
rect 377490 270444 377496 270456
rect 377548 270444 377554 270496
rect 378502 270444 378508 270496
rect 378560 270484 378566 270496
rect 379974 270484 379980 270496
rect 378560 270456 379980 270484
rect 378560 270444 378566 270456
rect 379974 270444 379980 270456
rect 380032 270444 380038 270496
rect 411254 270484 411260 270496
rect 380360 270456 411260 270484
rect 216916 270388 219434 270416
rect 216916 270376 216922 270388
rect 219894 270376 219900 270428
rect 219952 270416 219958 270428
rect 220262 270416 220268 270428
rect 219952 270388 220268 270416
rect 219952 270376 219958 270388
rect 220262 270376 220268 270388
rect 220320 270416 220326 270428
rect 245654 270416 245660 270428
rect 220320 270388 245660 270416
rect 220320 270376 220326 270388
rect 245654 270376 245660 270388
rect 245712 270376 245718 270428
rect 378042 270376 378048 270428
rect 378100 270416 378106 270428
rect 379238 270416 379244 270428
rect 378100 270388 379244 270416
rect 378100 270376 378106 270388
rect 379238 270376 379244 270388
rect 379296 270416 379302 270428
rect 380360 270416 380388 270456
rect 411254 270444 411260 270456
rect 411312 270444 411318 270496
rect 379296 270388 380388 270416
rect 379296 270376 379302 270388
rect 380434 270376 380440 270428
rect 380492 270416 380498 270428
rect 407114 270416 407120 270428
rect 380492 270388 407120 270416
rect 380492 270376 380498 270388
rect 407114 270376 407120 270388
rect 407172 270376 407178 270428
rect 51718 270308 51724 270360
rect 51776 270348 51782 270360
rect 84654 270348 84660 270360
rect 51776 270320 84660 270348
rect 51776 270308 51782 270320
rect 84654 270308 84660 270320
rect 84712 270308 84718 270360
rect 88242 270308 88248 270360
rect 88300 270348 88306 270360
rect 109034 270348 109040 270360
rect 88300 270320 109040 270348
rect 88300 270308 88306 270320
rect 109034 270308 109040 270320
rect 109092 270308 109098 270360
rect 217870 270308 217876 270360
rect 217928 270348 217934 270360
rect 249794 270348 249800 270360
rect 217928 270320 249800 270348
rect 217928 270308 217934 270320
rect 249794 270308 249800 270320
rect 249852 270308 249858 270360
rect 377950 270308 377956 270360
rect 378008 270348 378014 270360
rect 408494 270348 408500 270360
rect 378008 270320 408500 270348
rect 378008 270308 378014 270320
rect 408494 270308 408500 270320
rect 408552 270308 408558 270360
rect 59722 270240 59728 270292
rect 59780 270280 59786 270292
rect 61010 270280 61016 270292
rect 59780 270252 61016 270280
rect 59780 270240 59786 270252
rect 61010 270240 61016 270252
rect 61068 270240 61074 270292
rect 81434 270240 81440 270292
rect 81492 270280 81498 270292
rect 111794 270280 111800 270292
rect 81492 270252 111800 270280
rect 81492 270240 81498 270252
rect 111794 270240 111800 270252
rect 111852 270240 111858 270292
rect 213454 270240 213460 270292
rect 213512 270280 213518 270292
rect 244274 270280 244280 270292
rect 213512 270252 244280 270280
rect 213512 270240 213518 270252
rect 244274 270240 244280 270252
rect 244332 270240 244338 270292
rect 371602 270240 371608 270292
rect 371660 270280 371666 270292
rect 373166 270280 373172 270292
rect 371660 270252 373172 270280
rect 371660 270240 371666 270252
rect 373166 270240 373172 270252
rect 373224 270280 373230 270292
rect 400214 270280 400220 270292
rect 373224 270252 400220 270280
rect 373224 270240 373230 270252
rect 400214 270240 400220 270252
rect 400272 270240 400278 270292
rect 52730 270172 52736 270224
rect 52788 270212 52794 270224
rect 54570 270212 54576 270224
rect 52788 270184 54576 270212
rect 52788 270172 52794 270184
rect 54570 270172 54576 270184
rect 54628 270212 54634 270224
rect 85574 270212 85580 270224
rect 54628 270184 85580 270212
rect 54628 270172 54634 270184
rect 85574 270172 85580 270184
rect 85632 270172 85638 270224
rect 86862 270172 86868 270224
rect 86920 270212 86926 270224
rect 110414 270212 110420 270224
rect 86920 270184 110420 270212
rect 86920 270172 86926 270184
rect 110414 270172 110420 270184
rect 110472 270172 110478 270224
rect 220630 270172 220636 270224
rect 220688 270212 220694 270224
rect 248506 270212 248512 270224
rect 220688 270184 248512 270212
rect 220688 270172 220694 270184
rect 248506 270172 248512 270184
rect 248564 270172 248570 270224
rect 377030 270172 377036 270224
rect 377088 270212 377094 270224
rect 378594 270212 378600 270224
rect 377088 270184 378600 270212
rect 377088 270172 377094 270184
rect 378594 270172 378600 270184
rect 378652 270172 378658 270224
rect 378686 270172 378692 270224
rect 378744 270212 378750 270224
rect 401686 270212 401692 270224
rect 378744 270184 401692 270212
rect 378744 270172 378750 270184
rect 401686 270172 401692 270184
rect 401744 270172 401750 270224
rect 58618 270104 58624 270156
rect 58676 270144 58682 270156
rect 89714 270144 89720 270156
rect 58676 270116 89720 270144
rect 58676 270104 58682 270116
rect 89714 270104 89720 270116
rect 89772 270104 89778 270156
rect 210326 270104 210332 270156
rect 210384 270144 210390 270156
rect 213454 270144 213460 270156
rect 210384 270116 213460 270144
rect 210384 270104 210390 270116
rect 213454 270104 213460 270116
rect 213512 270104 213518 270156
rect 218422 270104 218428 270156
rect 218480 270144 218486 270156
rect 218606 270144 218612 270156
rect 218480 270116 218612 270144
rect 218480 270104 218486 270116
rect 218606 270104 218612 270116
rect 218664 270104 218670 270156
rect 220722 270104 220728 270156
rect 220780 270144 220786 270156
rect 251174 270144 251180 270156
rect 220780 270116 251180 270144
rect 220780 270104 220786 270116
rect 251174 270104 251180 270116
rect 251232 270104 251238 270156
rect 371050 270104 371056 270156
rect 371108 270144 371114 270156
rect 397454 270144 397460 270156
rect 371108 270116 378732 270144
rect 371108 270104 371114 270116
rect 59354 270036 59360 270088
rect 59412 270076 59418 270088
rect 92474 270076 92480 270088
rect 59412 270048 92480 270076
rect 59412 270036 59418 270048
rect 92474 270036 92480 270048
rect 92532 270036 92538 270088
rect 210234 270036 210240 270088
rect 210292 270076 210298 270088
rect 219710 270076 219716 270088
rect 210292 270048 219716 270076
rect 210292 270036 210298 270048
rect 219710 270036 219716 270048
rect 219768 270076 219774 270088
rect 252554 270076 252560 270088
rect 219768 270048 252560 270076
rect 219768 270036 219774 270048
rect 252554 270036 252560 270048
rect 252612 270036 252618 270088
rect 378704 270076 378732 270116
rect 378888 270116 397460 270144
rect 378888 270076 378916 270116
rect 397454 270104 397460 270116
rect 397512 270104 397518 270156
rect 378704 270048 378916 270076
rect 379606 270036 379612 270088
rect 379664 270076 379670 270088
rect 405734 270076 405740 270088
rect 379664 270048 405740 270076
rect 379664 270036 379670 270048
rect 405734 270036 405740 270048
rect 405792 270036 405798 270088
rect 54478 269968 54484 270020
rect 54536 270008 54542 270020
rect 55950 270008 55956 270020
rect 54536 269980 55956 270008
rect 54536 269968 54542 269980
rect 55950 269968 55956 269980
rect 56008 270008 56014 270020
rect 88334 270008 88340 270020
rect 56008 269980 88340 270008
rect 56008 269968 56014 269980
rect 88334 269968 88340 269980
rect 88392 269968 88398 270020
rect 217226 269968 217232 270020
rect 217284 270008 217290 270020
rect 218606 270008 218612 270020
rect 217284 269980 218612 270008
rect 217284 269968 217290 269980
rect 218606 269968 218612 269980
rect 218664 270008 218670 270020
rect 263594 270008 263600 270020
rect 218664 269980 263600 270008
rect 218664 269968 218670 269980
rect 263594 269968 263600 269980
rect 263652 269968 263658 270020
rect 374914 269968 374920 270020
rect 374972 270008 374978 270020
rect 379790 270008 379796 270020
rect 374972 269980 379796 270008
rect 374972 269968 374978 269980
rect 379790 269968 379796 269980
rect 379848 269968 379854 270020
rect 379974 269968 379980 270020
rect 380032 270008 380038 270020
rect 403618 270008 403624 270020
rect 380032 269980 403624 270008
rect 380032 269968 380038 269980
rect 403618 269968 403624 269980
rect 403676 269968 403682 270020
rect 80054 269900 80060 269952
rect 80112 269940 80118 269952
rect 114554 269940 114560 269952
rect 80112 269912 114560 269940
rect 80112 269900 80118 269912
rect 114554 269900 114560 269912
rect 114612 269900 114618 269952
rect 219342 269900 219348 269952
rect 219400 269940 219406 269952
rect 265158 269940 265164 269952
rect 219400 269912 265164 269940
rect 219400 269900 219406 269912
rect 265158 269900 265164 269912
rect 265216 269900 265222 269952
rect 368290 269900 368296 269952
rect 368348 269940 368354 269952
rect 398834 269940 398840 269952
rect 368348 269912 398840 269940
rect 368348 269900 368354 269912
rect 398834 269900 398840 269912
rect 398892 269900 398898 269952
rect 57238 269832 57244 269884
rect 57296 269872 57302 269884
rect 91094 269872 91100 269884
rect 57296 269844 91100 269872
rect 57296 269832 57302 269844
rect 91094 269832 91100 269844
rect 91152 269832 91158 269884
rect 113358 269832 113364 269884
rect 113416 269872 113422 269884
rect 128354 269872 128360 269884
rect 113416 269844 128360 269872
rect 113416 269832 113422 269844
rect 128354 269832 128360 269844
rect 128412 269832 128418 269884
rect 219066 269832 219072 269884
rect 219124 269872 219130 269884
rect 266354 269872 266360 269884
rect 219124 269844 266360 269872
rect 219124 269832 219130 269844
rect 266354 269832 266360 269844
rect 266412 269832 266418 269884
rect 378594 269832 378600 269884
rect 378652 269872 378658 269884
rect 411346 269872 411352 269884
rect 378652 269844 411352 269872
rect 378652 269832 378658 269844
rect 411346 269832 411352 269844
rect 411404 269832 411410 269884
rect 61010 269764 61016 269816
rect 61068 269804 61074 269816
rect 118694 269804 118700 269816
rect 61068 269776 118700 269804
rect 61068 269764 61074 269776
rect 118694 269764 118700 269776
rect 118752 269764 118758 269816
rect 213454 269764 213460 269816
rect 213512 269804 213518 269816
rect 271874 269804 271880 269816
rect 213512 269776 271880 269804
rect 213512 269764 213518 269776
rect 271874 269764 271880 269776
rect 271932 269764 271938 269816
rect 370958 269764 370964 269816
rect 371016 269804 371022 269816
rect 379974 269804 379980 269816
rect 371016 269776 379980 269804
rect 371016 269764 371022 269776
rect 379974 269764 379980 269776
rect 380032 269804 380038 269816
rect 413002 269804 413008 269816
rect 380032 269776 413008 269804
rect 380032 269764 380038 269776
rect 413002 269764 413008 269776
rect 413060 269764 413066 269816
rect 50614 269696 50620 269748
rect 50672 269736 50678 269748
rect 54662 269736 54668 269748
rect 50672 269708 54668 269736
rect 50672 269696 50678 269708
rect 54662 269696 54668 269708
rect 54720 269736 54726 269748
rect 84194 269736 84200 269748
rect 54720 269708 84200 269736
rect 54720 269696 54726 269708
rect 84194 269696 84200 269708
rect 84252 269696 84258 269748
rect 208210 269696 208216 269748
rect 208268 269736 208274 269748
rect 209406 269736 209412 269748
rect 208268 269708 209412 269736
rect 208268 269696 208274 269708
rect 209406 269696 209412 269708
rect 209464 269736 209470 269748
rect 237374 269736 237380 269748
rect 209464 269708 237380 269736
rect 209464 269696 209470 269708
rect 237374 269696 237380 269708
rect 237432 269696 237438 269748
rect 216582 269628 216588 269680
rect 216640 269668 216646 269680
rect 262214 269668 262220 269680
rect 216640 269640 262220 269668
rect 216640 269628 216646 269640
rect 262214 269628 262220 269640
rect 262272 269628 262278 269680
rect 219158 269560 219164 269612
rect 219216 269600 219222 269612
rect 219894 269600 219900 269612
rect 219216 269572 219900 269600
rect 219216 269560 219222 269572
rect 219894 269560 219900 269572
rect 219952 269600 219958 269612
rect 220722 269600 220728 269612
rect 219952 269572 220728 269600
rect 219952 269560 219958 269572
rect 220722 269560 220728 269572
rect 220780 269560 220786 269612
rect 251266 269600 251272 269612
rect 229066 269572 251272 269600
rect 218514 269492 218520 269544
rect 218572 269532 218578 269544
rect 219250 269532 219256 269544
rect 218572 269504 219256 269532
rect 218572 269492 218578 269504
rect 219250 269492 219256 269504
rect 219308 269532 219314 269544
rect 229066 269532 229094 269572
rect 251266 269560 251272 269572
rect 251324 269560 251330 269612
rect 375742 269560 375748 269612
rect 375800 269600 375806 269612
rect 376386 269600 376392 269612
rect 375800 269572 376392 269600
rect 375800 269560 375806 269572
rect 376386 269560 376392 269572
rect 376444 269600 376450 269612
rect 380434 269600 380440 269612
rect 376444 269572 380440 269600
rect 376444 269560 376450 269572
rect 380434 269560 380440 269572
rect 380492 269560 380498 269612
rect 219308 269504 229094 269532
rect 219308 269492 219314 269504
rect 218606 269356 218612 269408
rect 218664 269396 218670 269408
rect 219066 269396 219072 269408
rect 218664 269368 219072 269396
rect 218664 269356 218670 269368
rect 219066 269356 219072 269368
rect 219124 269356 219130 269408
rect 218146 269288 218152 269340
rect 218204 269328 218210 269340
rect 220262 269328 220268 269340
rect 218204 269300 220268 269328
rect 218204 269288 218210 269300
rect 220262 269288 220268 269300
rect 220320 269288 220326 269340
rect 214282 269220 214288 269272
rect 214340 269260 214346 269272
rect 219618 269260 219624 269272
rect 214340 269232 219624 269260
rect 214340 269220 214346 269232
rect 219618 269220 219624 269232
rect 219676 269260 219682 269272
rect 220630 269260 220636 269272
rect 219676 269232 220636 269260
rect 219676 269220 219682 269232
rect 220630 269220 220636 269232
rect 220688 269220 220694 269272
rect 375006 269192 375012 269204
rect 373966 269164 375012 269192
rect 219342 269084 219348 269136
rect 219400 269124 219406 269136
rect 219618 269124 219624 269136
rect 219400 269096 219624 269124
rect 219400 269084 219406 269096
rect 219618 269084 219624 269096
rect 219676 269084 219682 269136
rect 373626 269084 373632 269136
rect 373684 269124 373690 269136
rect 373966 269124 373994 269164
rect 375006 269152 375012 269164
rect 375064 269192 375070 269204
rect 378686 269192 378692 269204
rect 375064 269164 378692 269192
rect 375064 269152 375070 269164
rect 378686 269152 378692 269164
rect 378744 269152 378750 269204
rect 373684 269096 373994 269124
rect 373684 269084 373690 269096
rect 377490 269084 377496 269136
rect 377548 269124 377554 269136
rect 391934 269124 391940 269136
rect 377548 269096 391940 269124
rect 377548 269084 377554 269096
rect 391934 269084 391940 269096
rect 391992 269084 391998 269136
rect 47394 269016 47400 269068
rect 47452 269056 47458 269068
rect 58618 269056 58624 269068
rect 47452 269028 58624 269056
rect 47452 269016 47458 269028
rect 58618 269016 58624 269028
rect 58676 269016 58682 269068
rect 128354 269016 128360 269068
rect 128412 269056 128418 269068
rect 196986 269056 196992 269068
rect 128412 269028 196992 269056
rect 128412 269016 128418 269028
rect 196986 269016 196992 269028
rect 197044 269016 197050 269068
rect 208946 269016 208952 269068
rect 209004 269056 209010 269068
rect 217226 269056 217232 269068
rect 209004 269028 217232 269056
rect 209004 269016 209010 269028
rect 217226 269016 217232 269028
rect 217284 269056 217290 269068
rect 258074 269056 258080 269068
rect 217284 269028 258080 269056
rect 217284 269016 217290 269028
rect 258074 269016 258080 269028
rect 258132 269016 258138 269068
rect 375834 269016 375840 269068
rect 375892 269056 375898 269068
rect 416774 269056 416780 269068
rect 375892 269028 416780 269056
rect 375892 269016 375898 269028
rect 416774 269016 416780 269028
rect 416832 269016 416838 269068
rect 213638 268948 213644 269000
rect 213696 268988 213702 269000
rect 215846 268988 215852 269000
rect 213696 268960 215852 268988
rect 213696 268948 213702 268960
rect 215846 268948 215852 268960
rect 215904 268948 215910 269000
rect 216214 268948 216220 269000
rect 216272 268988 216278 269000
rect 216490 268988 216496 269000
rect 216272 268960 216496 268988
rect 216272 268948 216278 268960
rect 216490 268948 216496 268960
rect 216548 268948 216554 269000
rect 219434 268948 219440 269000
rect 219492 268988 219498 269000
rect 253934 268988 253940 269000
rect 219492 268960 253940 268988
rect 219492 268948 219498 268960
rect 253934 268948 253940 268960
rect 253992 268948 253998 269000
rect 375650 268948 375656 269000
rect 375708 268988 375714 269000
rect 375926 268988 375932 269000
rect 375708 268960 375932 268988
rect 375708 268948 375714 268960
rect 375926 268948 375932 268960
rect 375984 268948 375990 269000
rect 379882 268948 379888 269000
rect 379940 268988 379946 269000
rect 414014 268988 414020 269000
rect 379940 268960 414020 268988
rect 379940 268948 379946 268960
rect 414014 268948 414020 268960
rect 414072 268948 414078 269000
rect 216508 268920 216536 268948
rect 242894 268920 242900 268932
rect 216508 268892 242900 268920
rect 242894 268880 242900 268892
rect 242952 268880 242958 268932
rect 388438 268880 388444 268932
rect 388496 268920 388502 268932
rect 420914 268920 420920 268932
rect 388496 268892 420920 268920
rect 388496 268880 388502 268892
rect 420914 268880 420920 268892
rect 420972 268880 420978 268932
rect 214834 268812 214840 268864
rect 214892 268852 214898 268864
rect 218422 268852 218428 268864
rect 214892 268824 218428 268852
rect 214892 268812 214898 268824
rect 218422 268812 218428 268824
rect 218480 268852 218486 268864
rect 244366 268852 244372 268864
rect 218480 268824 244372 268852
rect 218480 268812 218486 268824
rect 244366 268812 244372 268824
rect 244424 268812 244430 268864
rect 379146 268812 379152 268864
rect 379204 268852 379210 268864
rect 409874 268852 409880 268864
rect 379204 268824 409880 268852
rect 379204 268812 379210 268824
rect 409874 268812 409880 268824
rect 409932 268812 409938 268864
rect 214374 268744 214380 268796
rect 214432 268784 214438 268796
rect 218514 268784 218520 268796
rect 214432 268756 218520 268784
rect 214432 268744 214438 268756
rect 218514 268744 218520 268756
rect 218572 268744 218578 268796
rect 235994 268784 236000 268796
rect 219406 268756 236000 268784
rect 215846 268676 215852 268728
rect 215904 268716 215910 268728
rect 219406 268716 219434 268756
rect 235994 268744 236000 268756
rect 236052 268744 236058 268796
rect 390554 268744 390560 268796
rect 390612 268784 390618 268796
rect 419534 268784 419540 268796
rect 390612 268756 419540 268784
rect 390612 268744 390618 268756
rect 419534 268744 419540 268756
rect 419592 268744 419598 268796
rect 215904 268688 219434 268716
rect 215904 268676 215910 268688
rect 232498 268676 232504 268728
rect 232556 268716 232562 268728
rect 259454 268716 259460 268728
rect 232556 268688 259460 268716
rect 232556 268676 232562 268688
rect 259454 268676 259460 268688
rect 259512 268676 259518 268728
rect 375926 268676 375932 268728
rect 375984 268716 375990 268728
rect 402974 268716 402980 268728
rect 375984 268688 402980 268716
rect 375984 268676 375990 268688
rect 402974 268676 402980 268688
rect 403032 268676 403038 268728
rect 43622 268608 43628 268660
rect 43680 268648 43686 268660
rect 46474 268648 46480 268660
rect 43680 268620 46480 268648
rect 43680 268608 43686 268620
rect 46474 268608 46480 268620
rect 46532 268648 46538 268660
rect 80054 268648 80060 268660
rect 46532 268620 80060 268648
rect 46532 268608 46538 268620
rect 80054 268608 80060 268620
rect 80112 268608 80118 268660
rect 213546 268608 213552 268660
rect 213604 268648 213610 268660
rect 217042 268648 217048 268660
rect 213604 268620 217048 268648
rect 213604 268608 213610 268620
rect 217042 268608 217048 268620
rect 217100 268608 217106 268660
rect 217410 268608 217416 268660
rect 217468 268648 217474 268660
rect 230474 268648 230480 268660
rect 217468 268620 230480 268648
rect 217468 268608 217474 268620
rect 230474 268608 230480 268620
rect 230532 268648 230538 268660
rect 259546 268648 259552 268660
rect 230532 268620 259552 268648
rect 230532 268608 230538 268620
rect 259546 268608 259552 268620
rect 259604 268608 259610 268660
rect 391934 268608 391940 268660
rect 391992 268648 391998 268660
rect 418154 268648 418160 268660
rect 391992 268620 418160 268648
rect 391992 268608 391998 268620
rect 418154 268608 418160 268620
rect 418212 268608 418218 268660
rect 43806 268540 43812 268592
rect 43864 268580 43870 268592
rect 46382 268580 46388 268592
rect 43864 268552 46388 268580
rect 43864 268540 43870 268552
rect 46382 268540 46388 268552
rect 46440 268580 46446 268592
rect 81434 268580 81440 268592
rect 46440 268552 81440 268580
rect 46440 268540 46446 268552
rect 81434 268540 81440 268552
rect 81492 268540 81498 268592
rect 229738 268540 229744 268592
rect 229796 268580 229802 268592
rect 260834 268580 260840 268592
rect 229796 268552 260840 268580
rect 229796 268540 229802 268552
rect 260834 268540 260840 268552
rect 260892 268540 260898 268592
rect 43530 268472 43536 268524
rect 43588 268512 43594 268524
rect 46198 268512 46204 268524
rect 43588 268484 46204 268512
rect 43588 268472 43594 268484
rect 46198 268472 46204 268484
rect 46256 268512 46262 268524
rect 86862 268512 86868 268524
rect 46256 268484 86868 268512
rect 46256 268472 46262 268484
rect 86862 268472 86868 268484
rect 86920 268472 86926 268524
rect 218514 268472 218520 268524
rect 218572 268512 218578 268524
rect 256694 268512 256700 268524
rect 218572 268484 256700 268512
rect 218572 268472 218578 268484
rect 256694 268472 256700 268484
rect 256752 268472 256758 268524
rect 43714 268404 43720 268456
rect 43772 268444 43778 268456
rect 46290 268444 46296 268456
rect 43772 268416 46296 268444
rect 43772 268404 43778 268416
rect 46290 268404 46296 268416
rect 46348 268444 46354 268456
rect 88242 268444 88248 268456
rect 46348 268416 88248 268444
rect 46348 268404 46354 268416
rect 88242 268404 88248 268416
rect 88300 268404 88306 268456
rect 217042 268404 217048 268456
rect 217100 268444 217106 268456
rect 255314 268444 255320 268456
rect 217100 268416 255320 268444
rect 217100 268404 217106 268416
rect 255314 268404 255320 268416
rect 255372 268404 255378 268456
rect 47578 268336 47584 268388
rect 47636 268376 47642 268388
rect 99374 268376 99380 268388
rect 47636 268348 99380 268376
rect 47636 268336 47642 268348
rect 99374 268336 99380 268348
rect 99432 268336 99438 268388
rect 202690 268336 202696 268388
rect 202748 268376 202754 268388
rect 212166 268376 212172 268388
rect 202748 268348 212172 268376
rect 202748 268336 202754 268348
rect 212166 268336 212172 268348
rect 212224 268376 212230 268388
rect 268194 268376 268200 268388
rect 212224 268348 268200 268376
rect 212224 268336 212230 268348
rect 268194 268336 268200 268348
rect 268252 268336 268258 268388
rect 372430 268336 372436 268388
rect 372488 268376 372494 268388
rect 374546 268376 374552 268388
rect 372488 268348 374552 268376
rect 372488 268336 372494 268348
rect 374546 268336 374552 268348
rect 374604 268376 374610 268388
rect 404354 268376 404360 268388
rect 374604 268348 404360 268376
rect 374604 268336 374610 268348
rect 404354 268336 404360 268348
rect 404412 268336 404418 268388
rect 43898 267656 43904 267708
rect 43956 267696 43962 267708
rect 47578 267696 47584 267708
rect 43956 267668 47584 267696
rect 43956 267656 43962 267668
rect 47578 267656 47584 267668
rect 47636 267656 47642 267708
rect 371694 267656 371700 267708
rect 371752 267696 371758 267708
rect 375190 267696 375196 267708
rect 371752 267668 375196 267696
rect 371752 267656 371758 267668
rect 375190 267656 375196 267668
rect 375248 267696 375254 267708
rect 434806 267696 434812 267708
rect 375248 267668 434812 267696
rect 375248 267656 375254 267668
rect 434806 267656 434812 267668
rect 434864 267656 434870 267708
rect 379054 267044 379060 267096
rect 379112 267084 379118 267096
rect 437474 267084 437480 267096
rect 379112 267056 437480 267084
rect 379112 267044 379118 267056
rect 437474 267044 437480 267056
rect 437532 267044 437538 267096
rect 373810 266976 373816 267028
rect 373868 267016 373874 267028
rect 375926 267016 375932 267028
rect 373868 266988 375932 267016
rect 373868 266976 373874 266988
rect 375926 266976 375932 266988
rect 375984 267016 375990 267028
rect 436094 267016 436100 267028
rect 375984 266988 436100 267016
rect 375984 266976 375990 266988
rect 436094 266976 436100 266988
rect 436152 266976 436158 267028
rect 219434 262896 219440 262948
rect 219492 262936 219498 262948
rect 219710 262936 219716 262948
rect 219492 262908 219716 262936
rect 219492 262896 219498 262908
rect 219710 262896 219716 262908
rect 219768 262896 219774 262948
rect 357066 253960 357072 253972
rect 356440 253932 357072 253960
rect 340782 253852 340788 253904
rect 340840 253892 340846 253904
rect 356440 253892 356468 253932
rect 357066 253920 357072 253932
rect 357124 253960 357130 253972
rect 357618 253960 357624 253972
rect 357124 253932 357624 253960
rect 357124 253920 357130 253932
rect 357618 253920 357624 253932
rect 357676 253920 357682 253972
rect 340840 253864 356468 253892
rect 340840 253852 340846 253864
rect 180150 253308 180156 253360
rect 180208 253348 180214 253360
rect 197538 253348 197544 253360
rect 180208 253320 197544 253348
rect 180208 253308 180214 253320
rect 197538 253308 197544 253320
rect 197596 253308 197602 253360
rect 500862 253308 500868 253360
rect 500920 253348 500926 253360
rect 517698 253348 517704 253360
rect 500920 253320 517704 253348
rect 500920 253308 500926 253320
rect 517698 253308 517704 253320
rect 517756 253308 517762 253360
rect 179322 253240 179328 253292
rect 179380 253280 179386 253292
rect 197354 253280 197360 253292
rect 179380 253252 197360 253280
rect 179380 253240 179386 253252
rect 197354 253240 197360 253252
rect 197412 253280 197418 253292
rect 197630 253280 197636 253292
rect 197412 253252 197636 253280
rect 197412 253240 197418 253252
rect 197630 253240 197636 253252
rect 197688 253240 197694 253292
rect 339402 253240 339408 253292
rect 339460 253280 339466 253292
rect 360194 253280 360200 253292
rect 339460 253252 360200 253280
rect 339460 253240 339466 253252
rect 360194 253240 360200 253252
rect 360252 253240 360258 253292
rect 499206 253240 499212 253292
rect 499264 253280 499270 253292
rect 517790 253280 517796 253292
rect 499264 253252 517796 253280
rect 499264 253240 499270 253252
rect 517790 253240 517796 253252
rect 517848 253240 517854 253292
rect 191742 253172 191748 253224
rect 191800 253212 191806 253224
rect 200758 253212 200764 253224
rect 191800 253184 200764 253212
rect 191800 253172 191806 253184
rect 200758 253172 200764 253184
rect 200816 253172 200822 253224
rect 351822 253172 351828 253224
rect 351880 253212 351886 253224
rect 358078 253212 358084 253224
rect 351880 253184 358084 253212
rect 351880 253172 351886 253184
rect 358078 253172 358084 253184
rect 358136 253172 358142 253224
rect 517698 253172 517704 253224
rect 517756 253212 517762 253224
rect 517974 253212 517980 253224
rect 517756 253184 517980 253212
rect 517756 253172 517762 253184
rect 517974 253172 517980 253184
rect 518032 253172 518038 253224
rect 510890 252560 510896 252612
rect 510948 252600 510954 252612
rect 517514 252600 517520 252612
rect 510948 252572 517520 252600
rect 510948 252560 510954 252572
rect 517514 252560 517520 252572
rect 517572 252560 517578 252612
rect 58802 252492 58808 252544
rect 58860 252532 58866 252544
rect 60918 252532 60924 252544
rect 58860 252504 60924 252532
rect 58860 252492 58866 252504
rect 60918 252492 60924 252504
rect 60976 252492 60982 252544
rect 214466 252492 214472 252544
rect 214524 252532 214530 252544
rect 214742 252532 214748 252544
rect 214524 252504 214748 252532
rect 214524 252492 214530 252504
rect 214742 252492 214748 252504
rect 214800 252492 214806 252544
rect 218606 252492 218612 252544
rect 218664 252532 218670 252544
rect 220814 252532 220820 252544
rect 218664 252504 220820 252532
rect 218664 252492 218670 252504
rect 220814 252492 220820 252504
rect 220872 252492 220878 252544
rect 232498 252532 232504 252544
rect 224236 252504 232504 252532
rect 56962 252424 56968 252476
rect 57020 252464 57026 252476
rect 61010 252464 61016 252476
rect 57020 252436 61016 252464
rect 57020 252424 57026 252436
rect 61010 252424 61016 252436
rect 61068 252424 61074 252476
rect 215754 252424 215760 252476
rect 215812 252464 215818 252476
rect 216398 252464 216404 252476
rect 215812 252436 216404 252464
rect 215812 252424 215818 252436
rect 216398 252424 216404 252436
rect 216456 252464 216462 252476
rect 224236 252464 224264 252504
rect 232498 252492 232504 252504
rect 232556 252492 232562 252544
rect 375282 252492 375288 252544
rect 375340 252532 375346 252544
rect 377398 252532 377404 252544
rect 375340 252504 377404 252532
rect 375340 252492 375346 252504
rect 377398 252492 377404 252504
rect 377456 252492 377462 252544
rect 378410 252492 378416 252544
rect 378468 252532 378474 252544
rect 434714 252532 434720 252544
rect 378468 252504 434720 252532
rect 378468 252492 378474 252504
rect 434714 252492 434720 252504
rect 434772 252492 434778 252544
rect 229738 252464 229744 252476
rect 216456 252436 224264 252464
rect 229066 252436 229744 252464
rect 216456 252424 216462 252436
rect 214742 252356 214748 252408
rect 214800 252396 214806 252408
rect 229066 252396 229094 252436
rect 229738 252424 229744 252436
rect 229796 252424 229802 252476
rect 371786 252424 371792 252476
rect 371844 252464 371850 252476
rect 373718 252464 373724 252476
rect 371844 252436 373724 252464
rect 371844 252424 371850 252436
rect 373718 252424 373724 252436
rect 373776 252464 373782 252476
rect 427078 252464 427084 252476
rect 373776 252436 427084 252464
rect 373776 252424 373782 252436
rect 427078 252424 427084 252436
rect 427136 252424 427142 252476
rect 214800 252368 229094 252396
rect 214800 252356 214806 252368
rect 375190 252356 375196 252408
rect 375248 252396 375254 252408
rect 376570 252396 376576 252408
rect 375248 252368 376576 252396
rect 375248 252356 375254 252368
rect 376570 252356 376576 252368
rect 376628 252356 376634 252408
rect 377398 252356 377404 252408
rect 377456 252396 377462 252408
rect 396718 252396 396724 252408
rect 377456 252368 396724 252396
rect 377456 252356 377462 252368
rect 396718 252356 396724 252368
rect 396776 252356 396782 252408
rect 376588 252328 376616 252356
rect 378410 252328 378416 252340
rect 376588 252300 378416 252328
rect 378410 252288 378416 252300
rect 378468 252288 378474 252340
rect 54478 251948 54484 252000
rect 54536 251988 54542 252000
rect 60734 251988 60740 252000
rect 54536 251960 60740 251988
rect 54536 251948 54542 251960
rect 60734 251948 60740 251960
rect 60792 251948 60798 252000
rect 58526 251880 58532 251932
rect 58584 251920 58590 251932
rect 106274 251920 106280 251932
rect 58584 251892 106280 251920
rect 58584 251880 58590 251892
rect 106274 251880 106280 251892
rect 106332 251880 106338 251932
rect 368382 251880 368388 251932
rect 368440 251920 368446 251932
rect 372246 251920 372252 251932
rect 368440 251892 372252 251920
rect 368440 251880 368446 251892
rect 372246 251880 372252 251892
rect 372304 251920 372310 251932
rect 425698 251920 425704 251932
rect 372304 251892 425704 251920
rect 372304 251880 372310 251892
rect 425698 251880 425704 251892
rect 425756 251880 425762 251932
rect 53834 251812 53840 251864
rect 53892 251852 53898 251864
rect 115934 251852 115940 251864
rect 53892 251824 115940 251852
rect 53892 251812 53898 251824
rect 115934 251812 115940 251824
rect 115992 251812 115998 251864
rect 216398 251812 216404 251864
rect 216456 251852 216462 251864
rect 230474 251852 230480 251864
rect 216456 251824 230480 251852
rect 216456 251812 216462 251824
rect 230474 251812 230480 251824
rect 230532 251812 230538 251864
rect 375282 251812 375288 251864
rect 375340 251852 375346 251864
rect 429194 251852 429200 251864
rect 375340 251824 429200 251852
rect 375340 251812 375346 251824
rect 429194 251812 429200 251824
rect 429252 251812 429258 251864
rect 58710 251608 58716 251660
rect 58768 251648 58774 251660
rect 60826 251648 60832 251660
rect 58768 251620 60832 251648
rect 58768 251608 58774 251620
rect 60826 251608 60832 251620
rect 60884 251608 60890 251660
rect 46842 251132 46848 251184
rect 46900 251172 46906 251184
rect 58526 251172 58532 251184
rect 46900 251144 58532 251172
rect 46900 251132 46906 251144
rect 58526 251132 58532 251144
rect 58584 251132 58590 251184
rect 372522 251132 372528 251184
rect 372580 251172 372586 251184
rect 374822 251172 374828 251184
rect 372580 251144 374828 251172
rect 372580 251132 372586 251144
rect 374822 251132 374828 251144
rect 374880 251172 374886 251184
rect 375282 251172 375288 251184
rect 374880 251144 375288 251172
rect 374880 251132 374886 251144
rect 375282 251132 375288 251144
rect 375340 251132 375346 251184
rect 49142 251064 49148 251116
rect 49200 251104 49206 251116
rect 53834 251104 53840 251116
rect 49200 251076 53840 251104
rect 49200 251064 49206 251076
rect 53834 251064 53840 251076
rect 53892 251104 53898 251116
rect 54294 251104 54300 251116
rect 53892 251076 54300 251104
rect 53892 251064 53898 251076
rect 54294 251064 54300 251076
rect 54352 251064 54358 251116
rect 519446 183540 519452 183592
rect 519504 183580 519510 183592
rect 520182 183580 520188 183592
rect 519504 183552 520188 183580
rect 519504 183540 519510 183552
rect 520182 183540 520188 183552
rect 520240 183580 520246 183592
rect 580258 183580 580264 183592
rect 520240 183552 580264 183580
rect 520240 183540 520246 183552
rect 580258 183540 580264 183552
rect 580316 183540 580322 183592
rect 520090 183472 520096 183524
rect 520148 183512 520154 183524
rect 580350 183512 580356 183524
rect 520148 183484 580356 183512
rect 520148 183472 520154 183484
rect 580350 183472 580356 183484
rect 580408 183472 580414 183524
rect 205082 177964 205088 178016
rect 205140 178004 205146 178016
rect 216674 178004 216680 178016
rect 205140 177976 216680 178004
rect 205140 177964 205146 177976
rect 216674 177964 216680 177976
rect 216732 177964 216738 178016
rect 365254 177964 365260 178016
rect 365312 178004 365318 178016
rect 376938 178004 376944 178016
rect 365312 177976 376944 178004
rect 365312 177964 365318 177976
rect 376938 177964 376944 177976
rect 376996 177964 377002 178016
rect 358078 175924 358084 175976
rect 358136 175964 358142 175976
rect 376938 175964 376944 175976
rect 358136 175936 376944 175964
rect 358136 175924 358142 175936
rect 376938 175924 376944 175936
rect 376996 175924 377002 175976
rect 216674 175284 216680 175296
rect 201512 175256 216680 175284
rect 201512 175228 201540 175256
rect 216674 175244 216680 175256
rect 216732 175244 216738 175296
rect 200758 175176 200764 175228
rect 200816 175216 200822 175228
rect 201494 175216 201500 175228
rect 200816 175188 201500 175216
rect 200816 175176 200822 175188
rect 201494 175176 201500 175188
rect 201552 175176 201558 175228
rect 207658 175176 207664 175228
rect 207716 175216 207722 175228
rect 216950 175216 216956 175228
rect 207716 175188 216956 175216
rect 207716 175176 207722 175188
rect 216950 175176 216956 175188
rect 217008 175176 217014 175228
rect 363782 175176 363788 175228
rect 363840 175216 363846 175228
rect 376938 175216 376944 175228
rect 363840 175188 376944 175216
rect 363840 175176 363846 175188
rect 376938 175176 376944 175188
rect 376996 175176 377002 175228
rect 50798 166948 50804 167000
rect 50856 166988 50862 167000
rect 96062 166988 96068 167000
rect 50856 166960 96068 166988
rect 50856 166948 50862 166960
rect 96062 166948 96068 166960
rect 96120 166948 96126 167000
rect 374638 166948 374644 167000
rect 374696 166988 374702 167000
rect 428274 166988 428280 167000
rect 374696 166960 428280 166988
rect 374696 166948 374702 166960
rect 428274 166948 428280 166960
rect 428332 166948 428338 167000
rect 49418 166880 49424 166932
rect 49476 166920 49482 166932
rect 98454 166920 98460 166932
rect 49476 166892 98460 166920
rect 49476 166880 49482 166892
rect 98454 166880 98460 166892
rect 98512 166880 98518 166932
rect 376202 166880 376208 166932
rect 376260 166920 376266 166932
rect 430942 166920 430948 166932
rect 376260 166892 430948 166920
rect 376260 166880 376266 166892
rect 430942 166880 430948 166892
rect 431000 166880 431006 166932
rect 50706 166812 50712 166864
rect 50764 166852 50770 166864
rect 101030 166852 101036 166864
rect 50764 166824 101036 166852
rect 50764 166812 50770 166824
rect 101030 166812 101036 166824
rect 101088 166812 101094 166864
rect 358354 166812 358360 166864
rect 358412 166852 358418 166864
rect 418430 166852 418436 166864
rect 358412 166824 418436 166852
rect 358412 166812 358418 166824
rect 418430 166812 418436 166824
rect 418488 166812 418494 166864
rect 53558 166744 53564 166796
rect 53616 166784 53622 166796
rect 105814 166784 105820 166796
rect 53616 166756 105820 166784
rect 53616 166744 53622 166756
rect 105814 166744 105820 166756
rect 105872 166744 105878 166796
rect 212166 166744 212172 166796
rect 212224 166784 212230 166796
rect 220814 166784 220820 166796
rect 212224 166756 220820 166784
rect 212224 166744 212230 166756
rect 220814 166744 220820 166756
rect 220872 166744 220878 166796
rect 358262 166744 358268 166796
rect 358320 166784 358326 166796
rect 421006 166784 421012 166796
rect 358320 166756 421012 166784
rect 358320 166744 358326 166756
rect 421006 166744 421012 166756
rect 421064 166744 421070 166796
rect 52178 166676 52184 166728
rect 52236 166716 52242 166728
rect 108206 166716 108212 166728
rect 52236 166688 108212 166716
rect 52236 166676 52242 166688
rect 108206 166676 108212 166688
rect 108264 166676 108270 166728
rect 210602 166676 210608 166728
rect 210660 166716 210666 166728
rect 260926 166716 260932 166728
rect 210660 166688 260932 166716
rect 210660 166676 210666 166688
rect 260926 166676 260932 166688
rect 260984 166676 260990 166728
rect 356698 166676 356704 166728
rect 356756 166716 356762 166728
rect 433610 166716 433616 166728
rect 356756 166688 433616 166716
rect 356756 166676 356762 166688
rect 433610 166676 433616 166688
rect 433668 166676 433674 166728
rect 59078 166608 59084 166660
rect 59136 166648 59142 166660
rect 140866 166648 140872 166660
rect 59136 166620 140872 166648
rect 59136 166608 59142 166620
rect 140866 166608 140872 166620
rect 140924 166608 140930 166660
rect 204898 166608 204904 166660
rect 204956 166648 204962 166660
rect 265894 166648 265900 166660
rect 204956 166620 265900 166648
rect 204956 166608 204962 166620
rect 265894 166608 265900 166620
rect 265952 166608 265958 166660
rect 372154 166608 372160 166660
rect 372212 166648 372218 166660
rect 475838 166648 475844 166660
rect 372212 166620 475844 166648
rect 372212 166608 372218 166620
rect 475838 166608 475844 166620
rect 475896 166608 475902 166660
rect 56226 166540 56232 166592
rect 56284 166580 56290 166592
rect 138474 166580 138480 166592
rect 56284 166552 138480 166580
rect 56284 166540 56290 166552
rect 138474 166540 138480 166552
rect 138532 166540 138538 166592
rect 204990 166540 204996 166592
rect 205048 166580 205054 166592
rect 288250 166580 288256 166592
rect 205048 166552 288256 166580
rect 205048 166540 205054 166552
rect 288250 166540 288256 166552
rect 288308 166540 288314 166592
rect 370682 166540 370688 166592
rect 370740 166580 370746 166592
rect 473446 166580 473452 166592
rect 370740 166552 473452 166580
rect 370740 166540 370746 166552
rect 473446 166540 473452 166552
rect 473504 166540 473510 166592
rect 59906 166472 59912 166524
rect 59964 166512 59970 166524
rect 145926 166512 145932 166524
rect 59964 166484 145932 166512
rect 59964 166472 59970 166484
rect 145926 166472 145932 166484
rect 145984 166472 145990 166524
rect 206462 166472 206468 166524
rect 206520 166512 206526 166524
rect 291010 166512 291016 166524
rect 206520 166484 291016 166512
rect 206520 166472 206526 166484
rect 291010 166472 291016 166484
rect 291068 166472 291074 166524
rect 373350 166472 373356 166524
rect 373408 166512 373414 166524
rect 480898 166512 480904 166524
rect 373408 166484 480904 166512
rect 373408 166472 373414 166484
rect 480898 166472 480904 166484
rect 480956 166472 480962 166524
rect 59170 166404 59176 166456
rect 59228 166444 59234 166456
rect 148502 166444 148508 166456
rect 59228 166416 148508 166444
rect 59228 166404 59234 166416
rect 148502 166404 148508 166416
rect 148560 166404 148566 166456
rect 202230 166404 202236 166456
rect 202288 166444 202294 166456
rect 285950 166444 285956 166456
rect 202288 166416 285956 166444
rect 202288 166404 202294 166416
rect 285950 166404 285956 166416
rect 286008 166404 286014 166456
rect 365162 166404 365168 166456
rect 365220 166444 365226 166456
rect 478414 166444 478420 166456
rect 365220 166416 478420 166444
rect 365220 166404 365226 166416
rect 478414 166404 478420 166416
rect 478472 166404 478478 166456
rect 58986 166336 58992 166388
rect 59044 166376 59050 166388
rect 153286 166376 153292 166388
rect 59044 166348 153292 166376
rect 59044 166336 59050 166348
rect 153286 166336 153292 166348
rect 153344 166336 153350 166388
rect 209130 166336 209136 166388
rect 209188 166376 209194 166388
rect 293310 166376 293316 166388
rect 209188 166348 293316 166376
rect 209188 166336 209194 166348
rect 293310 166336 293316 166348
rect 293368 166336 293374 166388
rect 367922 166336 367928 166388
rect 367980 166376 367986 166388
rect 483382 166376 483388 166388
rect 367980 166348 483388 166376
rect 367980 166336 367986 166348
rect 483382 166336 483388 166348
rect 483440 166336 483446 166388
rect 41322 166268 41328 166320
rect 41380 166308 41386 166320
rect 163314 166308 163320 166320
rect 41380 166280 163320 166308
rect 41380 166268 41386 166280
rect 163314 166268 163320 166280
rect 163372 166268 163378 166320
rect 211982 166268 211988 166320
rect 212040 166308 212046 166320
rect 298462 166308 298468 166320
rect 212040 166280 298468 166308
rect 212040 166268 212046 166280
rect 298462 166268 298468 166280
rect 298520 166268 298526 166320
rect 366634 166268 366640 166320
rect 366692 166308 366698 166320
rect 485958 166308 485964 166320
rect 366692 166280 485964 166308
rect 366692 166268 366698 166280
rect 485958 166268 485964 166280
rect 486016 166268 486022 166320
rect 54386 166200 54392 166252
rect 54444 166240 54450 166252
rect 60734 166240 60740 166252
rect 54444 166212 60740 166240
rect 54444 166200 54450 166212
rect 60734 166200 60740 166212
rect 60792 166200 60798 166252
rect 369394 166200 369400 166252
rect 369452 166240 369458 166252
rect 423398 166240 423404 166252
rect 369452 166212 423404 166240
rect 369452 166200 369458 166212
rect 423398 166200 423404 166212
rect 423456 166200 423462 166252
rect 357250 165792 357256 165844
rect 357308 165832 357314 165844
rect 360286 165832 360292 165844
rect 357308 165804 360292 165832
rect 357308 165792 357314 165804
rect 360286 165792 360292 165804
rect 360344 165792 360350 165844
rect 46198 165656 46204 165708
rect 46256 165696 46262 165708
rect 52178 165696 52184 165708
rect 46256 165668 52184 165696
rect 46256 165656 46262 165668
rect 52178 165656 52184 165668
rect 52236 165696 52242 165708
rect 111150 165696 111156 165708
rect 52236 165668 111156 165696
rect 52236 165656 52242 165668
rect 111150 165656 111156 165668
rect 111208 165656 111214 165708
rect 54294 165588 54300 165640
rect 54352 165628 54358 165640
rect 116946 165628 116952 165640
rect 54352 165600 116952 165628
rect 54352 165588 54358 165600
rect 116946 165588 116952 165600
rect 117004 165588 117010 165640
rect 356974 165628 356980 165640
rect 356348 165600 356980 165628
rect 59814 165520 59820 165572
rect 59872 165560 59878 165572
rect 150434 165560 150440 165572
rect 59872 165532 150440 165560
rect 59872 165520 59878 165532
rect 150434 165520 150440 165532
rect 150492 165520 150498 165572
rect 197354 165520 197360 165572
rect 197412 165560 197418 165572
rect 197722 165560 197728 165572
rect 197412 165532 197728 165560
rect 197412 165520 197418 165532
rect 197722 165520 197728 165532
rect 197780 165520 197786 165572
rect 216030 165520 216036 165572
rect 216088 165560 216094 165572
rect 325878 165560 325884 165572
rect 216088 165532 325884 165560
rect 216088 165520 216094 165532
rect 325878 165520 325884 165532
rect 325936 165520 325942 165572
rect 343266 165520 343272 165572
rect 343324 165560 343330 165572
rect 356348 165560 356376 165600
rect 356974 165588 356980 165600
rect 357032 165628 357038 165640
rect 357526 165628 357532 165640
rect 357032 165600 357532 165628
rect 357032 165588 357038 165600
rect 357526 165588 357532 165600
rect 357584 165588 357590 165640
rect 375282 165588 375288 165640
rect 375340 165628 375346 165640
rect 434346 165628 434352 165640
rect 375340 165600 434352 165628
rect 375340 165588 375346 165600
rect 434346 165588 434352 165600
rect 434404 165588 434410 165640
rect 343324 165532 356376 165560
rect 343324 165520 343330 165532
rect 362402 165520 362408 165572
rect 362460 165560 362466 165572
rect 458358 165560 458364 165572
rect 362460 165532 458364 165560
rect 362460 165520 362466 165532
rect 458358 165520 458364 165532
rect 458416 165520 458422 165572
rect 56134 165452 56140 165504
rect 56192 165492 56198 165504
rect 135254 165492 135260 165504
rect 56192 165464 135260 165492
rect 56192 165452 56198 165464
rect 135254 165452 135260 165464
rect 135312 165452 135318 165504
rect 210510 165452 210516 165504
rect 210568 165492 210574 165504
rect 320910 165492 320916 165504
rect 210568 165464 320916 165492
rect 210568 165452 210574 165464
rect 320910 165452 320916 165464
rect 320968 165452 320974 165504
rect 360930 165452 360936 165504
rect 360988 165492 360994 165504
rect 452654 165492 452660 165504
rect 360988 165464 452660 165492
rect 360988 165452 360994 165464
rect 452654 165452 452660 165464
rect 452712 165452 452718 165504
rect 55122 165384 55128 165436
rect 55180 165424 55186 165436
rect 132494 165424 132500 165436
rect 55180 165396 132500 165424
rect 55180 165384 55186 165396
rect 132494 165384 132500 165396
rect 132552 165384 132558 165436
rect 213178 165384 213184 165436
rect 213236 165424 213242 165436
rect 300854 165424 300860 165436
rect 213236 165396 300860 165424
rect 213236 165384 213242 165396
rect 300854 165384 300860 165396
rect 300912 165384 300918 165436
rect 369210 165384 369216 165436
rect 369268 165424 369274 165436
rect 455414 165424 455420 165436
rect 369268 165396 455420 165424
rect 369268 165384 369274 165396
rect 455414 165384 455420 165396
rect 455472 165384 455478 165436
rect 54846 165316 54852 165368
rect 54904 165356 54910 165368
rect 128354 165356 128360 165368
rect 54904 165328 128360 165356
rect 54904 165316 54910 165328
rect 128354 165316 128360 165328
rect 128412 165316 128418 165368
rect 214650 165316 214656 165368
rect 214708 165356 214714 165368
rect 280154 165356 280160 165368
rect 214708 165328 280160 165356
rect 214708 165316 214714 165328
rect 280154 165316 280160 165328
rect 280212 165316 280218 165368
rect 363690 165316 363696 165368
rect 363748 165356 363754 165368
rect 443454 165356 443460 165368
rect 363748 165328 443460 165356
rect 363748 165316 363754 165328
rect 443454 165316 443460 165328
rect 443512 165316 443518 165368
rect 56502 165248 56508 165300
rect 56560 165288 56566 165300
rect 129734 165288 129740 165300
rect 56560 165260 129740 165288
rect 56560 165248 56566 165260
rect 129734 165248 129740 165260
rect 129792 165248 129798 165300
rect 211890 165248 211896 165300
rect 211948 165288 211954 165300
rect 277394 165288 277400 165300
rect 211948 165260 277400 165288
rect 211948 165248 211954 165260
rect 277394 165248 277400 165260
rect 277452 165248 277458 165300
rect 370590 165248 370596 165300
rect 370648 165288 370654 165300
rect 449894 165288 449900 165300
rect 370648 165260 449900 165288
rect 370648 165248 370654 165260
rect 449894 165248 449900 165260
rect 449952 165248 449958 165300
rect 56318 165180 56324 165232
rect 56376 165220 56382 165232
rect 125870 165220 125876 165232
rect 56376 165192 125876 165220
rect 56376 165180 56382 165192
rect 125870 165180 125876 165192
rect 125928 165180 125934 165232
rect 218974 165180 218980 165232
rect 219032 165220 219038 165232
rect 283374 165220 283380 165232
rect 219032 165192 283380 165220
rect 219032 165180 219038 165192
rect 283374 165180 283380 165192
rect 283432 165180 283438 165232
rect 372062 165180 372068 165232
rect 372120 165220 372126 165232
rect 447318 165220 447324 165232
rect 372120 165192 447324 165220
rect 372120 165180 372126 165192
rect 447318 165180 447324 165192
rect 447376 165180 447382 165232
rect 55030 165112 55036 165164
rect 55088 165152 55094 165164
rect 123478 165152 123484 165164
rect 55088 165124 123484 165152
rect 55088 165112 55094 165124
rect 123478 165112 123484 165124
rect 123536 165112 123542 165164
rect 183462 165112 183468 165164
rect 183520 165152 183526 165164
rect 197354 165152 197360 165164
rect 183520 165124 197360 165152
rect 183520 165112 183526 165124
rect 197354 165112 197360 165124
rect 197412 165112 197418 165164
rect 206370 165112 206376 165164
rect 206428 165152 206434 165164
rect 267734 165152 267740 165164
rect 206428 165124 267740 165152
rect 206428 165112 206434 165124
rect 267734 165112 267740 165124
rect 267792 165112 267798 165164
rect 373258 165112 373264 165164
rect 373316 165152 373322 165164
rect 445846 165152 445852 165164
rect 373316 165124 445852 165152
rect 373316 165112 373322 165124
rect 445846 165112 445852 165124
rect 445904 165112 445910 165164
rect 503254 165112 503260 165164
rect 503312 165152 503318 165164
rect 517606 165152 517612 165164
rect 503312 165124 517612 165152
rect 503312 165112 503318 165124
rect 517606 165112 517612 165124
rect 517664 165112 517670 165164
rect 56042 165044 56048 165096
rect 56100 165084 56106 165096
rect 120902 165084 120908 165096
rect 56100 165056 120908 165084
rect 56100 165044 56106 165056
rect 120902 165044 120908 165056
rect 120960 165044 120966 165096
rect 218882 165044 218888 165096
rect 218940 165084 218946 165096
rect 276014 165084 276020 165096
rect 218940 165056 276020 165084
rect 218940 165044 218946 165056
rect 276014 165044 276020 165056
rect 276072 165044 276078 165096
rect 366542 165044 366548 165096
rect 366600 165084 366606 165096
rect 438486 165084 438492 165096
rect 366600 165056 438492 165084
rect 366600 165044 366606 165056
rect 438486 165044 438492 165056
rect 438544 165044 438550 165096
rect 440142 165044 440148 165096
rect 440200 165084 440206 165096
rect 516594 165084 516600 165096
rect 440200 165056 516600 165084
rect 440200 165044 440206 165056
rect 516594 165044 516600 165056
rect 516652 165044 516658 165096
rect 52086 164976 52092 165028
rect 52144 165016 52150 165028
rect 115934 165016 115940 165028
rect 52144 164988 115940 165016
rect 52144 164976 52150 164988
rect 115934 164976 115940 164988
rect 115992 164976 115998 165028
rect 183186 164976 183192 165028
rect 183244 165016 183250 165028
rect 197446 165016 197452 165028
rect 183244 164988 197452 165016
rect 183244 164976 183250 164988
rect 197446 164976 197452 164988
rect 197504 164976 197510 165028
rect 216122 164976 216128 165028
rect 216180 165016 216186 165028
rect 273438 165016 273444 165028
rect 216180 164988 273444 165016
rect 216180 164976 216186 164988
rect 273438 164976 273444 164988
rect 273496 164976 273502 165028
rect 367830 164976 367836 165028
rect 367888 165016 367894 165028
rect 435910 165016 435916 165028
rect 367888 164988 435916 165016
rect 367888 164976 367894 164988
rect 435910 164976 435916 164988
rect 435968 164976 435974 165028
rect 503346 164976 503352 165028
rect 503404 165016 503410 165028
rect 517882 165016 517888 165028
rect 503404 164988 517888 165016
rect 503404 164976 503410 164988
rect 517882 164976 517888 164988
rect 517940 164976 517946 165028
rect 54938 164908 54944 164960
rect 54996 164948 55002 164960
rect 113542 164948 113548 164960
rect 54996 164920 113548 164948
rect 54996 164908 55002 164920
rect 113542 164908 113548 164920
rect 113600 164908 113606 164960
rect 114646 164908 114652 164960
rect 114704 164948 114710 164960
rect 196710 164948 196716 164960
rect 114704 164920 196716 164948
rect 114704 164908 114710 164920
rect 196710 164908 196716 164920
rect 196768 164908 196774 164960
rect 202322 164908 202328 164960
rect 202380 164948 202386 164960
rect 255314 164948 255320 164960
rect 202380 164920 255320 164948
rect 202380 164908 202386 164920
rect 255314 164908 255320 164920
rect 255372 164908 255378 164960
rect 374730 164908 374736 164960
rect 374788 164948 374794 164960
rect 440878 164948 440884 164960
rect 374788 164920 440884 164948
rect 374788 164908 374794 164920
rect 440878 164908 440884 164920
rect 440936 164908 440942 164960
rect 510522 164908 510528 164960
rect 510580 164948 510586 164960
rect 517514 164948 517520 164960
rect 510580 164920 517520 164948
rect 510580 164908 510586 164920
rect 517514 164908 517520 164920
rect 517572 164908 517578 164960
rect 51994 164840 52000 164892
rect 52052 164880 52058 164892
rect 91738 164880 91744 164892
rect 52052 164852 91744 164880
rect 52052 164840 52058 164852
rect 91738 164840 91744 164852
rect 91796 164840 91802 164892
rect 114462 164840 114468 164892
rect 114520 164880 114526 164892
rect 114738 164880 114744 164892
rect 114520 164852 114744 164880
rect 114520 164840 114526 164852
rect 114738 164840 114744 164852
rect 114796 164880 114802 164892
rect 196618 164880 196624 164892
rect 114796 164852 196624 164880
rect 114796 164840 114802 164852
rect 196618 164840 196624 164852
rect 196676 164840 196682 164892
rect 203518 164840 203524 164892
rect 203576 164880 203582 164892
rect 249794 164880 249800 164892
rect 203576 164852 249800 164880
rect 203576 164840 203582 164852
rect 249794 164840 249800 164852
rect 249852 164840 249858 164892
rect 343450 164840 343456 164892
rect 343508 164880 343514 164892
rect 356698 164880 356704 164892
rect 343508 164852 356704 164880
rect 343508 164840 343514 164852
rect 356698 164840 356704 164852
rect 356756 164880 356762 164892
rect 357250 164880 357256 164892
rect 356756 164852 357256 164880
rect 356756 164840 356762 164852
rect 357250 164840 357256 164852
rect 357308 164840 357314 164892
rect 365070 164840 365076 164892
rect 365128 164880 365134 164892
rect 412634 164880 412640 164892
rect 365128 164852 412640 164880
rect 365128 164840 365134 164852
rect 412634 164840 412640 164852
rect 412692 164840 412698 164892
rect 53466 164772 53472 164824
rect 53524 164812 53530 164824
rect 94590 164812 94596 164824
rect 53524 164784 94596 164812
rect 53524 164772 53530 164784
rect 94590 164772 94596 164784
rect 94648 164772 94654 164824
rect 94774 164772 94780 164824
rect 94832 164812 94838 164824
rect 118142 164812 118148 164824
rect 94832 164784 118148 164812
rect 94832 164772 94838 164784
rect 118142 164772 118148 164784
rect 118200 164772 118206 164824
rect 215938 164772 215944 164824
rect 215996 164812 216002 164824
rect 258074 164812 258080 164824
rect 215996 164784 258080 164812
rect 215996 164772 216002 164784
rect 258074 164772 258080 164784
rect 258132 164772 258138 164824
rect 378870 164772 378876 164824
rect 378928 164812 378934 164824
rect 416038 164812 416044 164824
rect 378928 164784 416044 164812
rect 378928 164772 378934 164784
rect 416038 164772 416044 164784
rect 416096 164772 416102 164824
rect 50890 164704 50896 164756
rect 50948 164744 50954 164756
rect 89990 164744 89996 164756
rect 50948 164716 89996 164744
rect 50948 164704 50954 164716
rect 89990 164704 89996 164716
rect 90048 164704 90054 164756
rect 211798 164704 211804 164756
rect 211856 164744 211862 164756
rect 252554 164744 252560 164756
rect 211856 164716 252560 164744
rect 211856 164704 211862 164716
rect 252554 164704 252560 164716
rect 252612 164704 252618 164756
rect 376110 164704 376116 164756
rect 376168 164744 376174 164756
rect 409874 164744 409880 164756
rect 376168 164716 409880 164744
rect 376168 164704 376174 164716
rect 409874 164704 409880 164716
rect 409932 164704 409938 164756
rect 56410 164636 56416 164688
rect 56468 164676 56474 164688
rect 88334 164676 88340 164688
rect 56468 164648 88340 164676
rect 56468 164636 56474 164648
rect 88334 164636 88340 164648
rect 88392 164636 88398 164688
rect 91738 164636 91744 164688
rect 91796 164676 91802 164688
rect 103514 164676 103520 164688
rect 91796 164648 103520 164676
rect 91796 164636 91802 164648
rect 103514 164636 103520 164648
rect 103572 164636 103578 164688
rect 214558 164636 214564 164688
rect 214616 164676 214622 164688
rect 247034 164676 247040 164688
rect 214616 164648 247040 164676
rect 214616 164636 214622 164648
rect 247034 164636 247040 164648
rect 247092 164636 247098 164688
rect 378962 164636 378968 164688
rect 379020 164676 379026 164688
rect 407114 164676 407120 164688
rect 379020 164648 407120 164676
rect 379020 164636 379026 164648
rect 407114 164636 407120 164648
rect 407172 164636 407178 164688
rect 98638 164296 98644 164348
rect 98696 164336 98702 164348
rect 100754 164336 100760 164348
rect 98696 164308 100760 164336
rect 98696 164296 98702 164308
rect 100754 164296 100760 164308
rect 100812 164296 100818 164348
rect 427814 164296 427820 164348
rect 427872 164336 427878 164348
rect 435082 164336 435088 164348
rect 427872 164308 435088 164336
rect 427872 164296 427878 164308
rect 435082 164296 435088 164308
rect 435140 164296 435146 164348
rect 100018 164228 100024 164280
rect 100076 164268 100082 164280
rect 103514 164268 103520 164280
rect 100076 164240 103520 164268
rect 100076 164228 100082 164240
rect 103514 164228 103520 164240
rect 103572 164228 103578 164280
rect 58526 164160 58532 164212
rect 58584 164200 58590 164212
rect 59906 164200 59912 164212
rect 58584 164172 59912 164200
rect 58584 164160 58590 164172
rect 59906 164160 59912 164172
rect 59964 164160 59970 164212
rect 117866 164200 117872 164212
rect 60016 164172 117872 164200
rect 57514 164092 57520 164144
rect 57572 164132 57578 164144
rect 60016 164132 60044 164172
rect 117866 164160 117872 164172
rect 117924 164160 117930 164212
rect 219618 164160 219624 164212
rect 219676 164200 219682 164212
rect 264974 164200 264980 164212
rect 219676 164172 264980 164200
rect 219676 164160 219682 164172
rect 264974 164160 264980 164172
rect 265032 164160 265038 164212
rect 374822 164160 374828 164212
rect 374880 164200 374886 164212
rect 429654 164200 429660 164212
rect 374880 164172 429660 164200
rect 374880 164160 374886 164172
rect 429654 164160 429660 164172
rect 429712 164160 429718 164212
rect 110966 164132 110972 164144
rect 57572 164104 60044 164132
rect 64846 164104 110972 164132
rect 57572 164092 57578 164104
rect 56962 163956 56968 164008
rect 57020 163996 57026 164008
rect 59446 163996 59452 164008
rect 57020 163968 59452 163996
rect 57020 163956 57026 163968
rect 59446 163956 59452 163968
rect 59504 163956 59510 164008
rect 53650 163888 53656 163940
rect 53708 163928 53714 163940
rect 64846 163928 64874 164104
rect 110966 164092 110972 164104
rect 111024 164092 111030 164144
rect 218330 164092 218336 164144
rect 218388 164132 218394 164144
rect 219066 164132 219072 164144
rect 218388 164104 219072 164132
rect 218388 164092 218394 164104
rect 219066 164092 219072 164104
rect 219124 164132 219130 164144
rect 263778 164132 263784 164144
rect 219124 164104 263784 164132
rect 219124 164092 219130 164104
rect 263778 164092 263784 164104
rect 263836 164092 263842 164144
rect 374454 164092 374460 164144
rect 374512 164132 374518 164144
rect 376110 164132 376116 164144
rect 374512 164104 376116 164132
rect 374512 164092 374518 164104
rect 376110 164092 376116 164104
rect 376168 164092 376174 164144
rect 379698 164092 379704 164144
rect 379756 164132 379762 164144
rect 426434 164132 426440 164144
rect 379756 164104 426440 164132
rect 379756 164092 379762 164104
rect 426434 164092 426440 164104
rect 426492 164092 426498 164144
rect 213362 164024 213368 164076
rect 213420 164064 213426 164076
rect 236086 164064 236092 164076
rect 213420 164036 236092 164064
rect 213420 164024 213426 164036
rect 236086 164024 236092 164036
rect 236144 164024 236150 164076
rect 379514 164024 379520 164076
rect 379572 164064 379578 164076
rect 426526 164064 426532 164076
rect 379572 164036 426532 164064
rect 379572 164024 379578 164036
rect 426526 164024 426532 164036
rect 426584 164024 426590 164076
rect 374914 163956 374920 164008
rect 374972 163996 374978 164008
rect 396166 163996 396172 164008
rect 374972 163968 396172 163996
rect 374972 163956 374978 163968
rect 396166 163956 396172 163968
rect 396224 163956 396230 164008
rect 53708 163900 64874 163928
rect 53708 163888 53714 163900
rect 212258 163888 212264 163940
rect 212316 163928 212322 163940
rect 213362 163928 213368 163940
rect 212316 163900 213368 163928
rect 212316 163888 212322 163900
rect 213362 163888 213368 163900
rect 213420 163888 213426 163940
rect 374362 163888 374368 163940
rect 374420 163928 374426 163940
rect 396074 163928 396080 163940
rect 374420 163900 396080 163928
rect 374420 163888 374426 163900
rect 396074 163888 396080 163900
rect 396132 163888 396138 163940
rect 51442 163820 51448 163872
rect 51500 163860 51506 163872
rect 57054 163860 57060 163872
rect 51500 163832 57060 163860
rect 51500 163820 51506 163832
rect 57054 163820 57060 163832
rect 57112 163860 57118 163872
rect 95234 163860 95240 163872
rect 57112 163832 95240 163860
rect 57112 163820 57118 163832
rect 95234 163820 95240 163832
rect 95292 163820 95298 163872
rect 50154 163752 50160 163804
rect 50212 163792 50218 163804
rect 56502 163792 56508 163804
rect 50212 163764 56508 163792
rect 50212 163752 50218 163764
rect 56502 163752 56508 163764
rect 56560 163792 56566 163804
rect 96614 163792 96620 163804
rect 56560 163764 96620 163792
rect 56560 163752 56566 163764
rect 96614 163752 96620 163764
rect 96672 163752 96678 163804
rect 48958 163684 48964 163736
rect 49016 163724 49022 163736
rect 55030 163724 55036 163736
rect 49016 163696 55036 163724
rect 49016 163684 49022 163696
rect 55030 163684 55036 163696
rect 55088 163724 55094 163736
rect 97994 163724 98000 163736
rect 55088 163696 98000 163724
rect 55088 163684 55094 163696
rect 97994 163684 98000 163696
rect 98052 163684 98058 163736
rect 59906 163616 59912 163668
rect 59964 163656 59970 163668
rect 106366 163656 106372 163668
rect 59964 163628 106372 163656
rect 59964 163616 59970 163628
rect 106366 163616 106372 163628
rect 106424 163616 106430 163668
rect 46290 163548 46296 163600
rect 46348 163588 46354 163600
rect 53650 163588 53656 163600
rect 46348 163560 53656 163588
rect 46348 163548 46354 163560
rect 53650 163548 53656 163560
rect 53708 163588 53714 163600
rect 109310 163588 109316 163600
rect 53708 163560 109316 163588
rect 53708 163548 53714 163560
rect 109310 163548 109316 163560
rect 109368 163548 109374 163600
rect 376110 163548 376116 163600
rect 376168 163588 376174 163600
rect 422294 163588 422300 163600
rect 376168 163560 422300 163588
rect 376168 163548 376174 163560
rect 422294 163548 422300 163560
rect 422352 163548 422358 163600
rect 59446 163480 59452 163532
rect 59504 163520 59510 163532
rect 118878 163520 118884 163532
rect 59504 163492 118884 163520
rect 59504 163480 59510 163492
rect 118878 163480 118884 163492
rect 118936 163480 118942 163532
rect 213362 163480 213368 163532
rect 213420 163520 213426 163532
rect 273806 163520 273812 163532
rect 213420 163492 273812 163520
rect 213420 163480 213426 163492
rect 273806 163480 273812 163492
rect 273864 163480 273870 163532
rect 371786 163480 371792 163532
rect 371844 163520 371850 163532
rect 374914 163520 374920 163532
rect 371844 163492 374920 163520
rect 371844 163480 371850 163492
rect 374914 163480 374920 163492
rect 374972 163520 374978 163532
rect 432230 163520 432236 163532
rect 374972 163492 432236 163520
rect 374972 163480 374978 163492
rect 432230 163480 432236 163492
rect 432288 163480 432294 163532
rect 46474 162800 46480 162852
rect 46532 162840 46538 162852
rect 50890 162840 50896 162852
rect 46532 162812 50896 162840
rect 46532 162800 46538 162812
rect 50890 162800 50896 162812
rect 50948 162800 50954 162852
rect 217042 162800 217048 162852
rect 217100 162840 217106 162852
rect 217870 162840 217876 162852
rect 217100 162812 217876 162840
rect 217100 162800 217106 162812
rect 217870 162800 217876 162812
rect 217928 162800 217934 162852
rect 218514 162800 218520 162852
rect 218572 162840 218578 162852
rect 218974 162840 218980 162852
rect 218572 162812 218980 162840
rect 218572 162800 218578 162812
rect 218974 162800 218980 162812
rect 219032 162800 219038 162852
rect 260834 162840 260840 162852
rect 219084 162812 260840 162840
rect 46382 162732 46388 162784
rect 46440 162772 46446 162784
rect 52086 162772 52092 162784
rect 46440 162744 52092 162772
rect 46440 162732 46446 162744
rect 52086 162732 52092 162744
rect 52144 162732 52150 162784
rect 214742 162732 214748 162784
rect 214800 162772 214806 162784
rect 219084 162772 219112 162812
rect 260834 162800 260840 162812
rect 260892 162800 260898 162852
rect 371694 162800 371700 162852
rect 371752 162840 371758 162852
rect 372522 162840 372528 162852
rect 371752 162812 372528 162840
rect 371752 162800 371758 162812
rect 372522 162800 372528 162812
rect 372580 162800 372586 162852
rect 375926 162800 375932 162852
rect 375984 162840 375990 162852
rect 376570 162840 376576 162852
rect 375984 162812 376576 162840
rect 375984 162800 375990 162812
rect 376570 162800 376576 162812
rect 376628 162800 376634 162852
rect 377490 162800 377496 162852
rect 377548 162840 377554 162852
rect 379606 162840 379612 162852
rect 377548 162812 379612 162840
rect 377548 162800 377554 162812
rect 379606 162800 379612 162812
rect 379664 162800 379670 162852
rect 379790 162800 379796 162852
rect 379848 162840 379854 162852
rect 436186 162840 436192 162852
rect 379848 162812 436192 162840
rect 379848 162800 379854 162812
rect 436186 162800 436192 162812
rect 436244 162800 436250 162852
rect 214800 162744 219112 162772
rect 214800 162732 214806 162744
rect 219342 162732 219348 162784
rect 219400 162772 219406 162784
rect 259454 162772 259460 162784
rect 219400 162744 259460 162772
rect 219400 162732 219406 162744
rect 259454 162732 259460 162744
rect 259512 162732 259518 162784
rect 375834 162732 375840 162784
rect 375892 162772 375898 162784
rect 378962 162772 378968 162784
rect 375892 162744 378968 162772
rect 375892 162732 375898 162744
rect 378962 162732 378968 162744
rect 379020 162732 379026 162784
rect 379054 162732 379060 162784
rect 379112 162772 379118 162784
rect 437934 162772 437940 162784
rect 379112 162744 437940 162772
rect 379112 162732 379118 162744
rect 437934 162732 437940 162744
rect 437992 162732 437998 162784
rect 216398 162664 216404 162716
rect 216456 162704 216462 162716
rect 259546 162704 259552 162716
rect 216456 162676 259552 162704
rect 216456 162664 216462 162676
rect 259546 162664 259552 162676
rect 259604 162664 259610 162716
rect 372522 162664 372528 162716
rect 372580 162704 372586 162716
rect 427814 162704 427820 162716
rect 372580 162676 427820 162704
rect 372580 162664 372586 162676
rect 427814 162664 427820 162676
rect 427872 162664 427878 162716
rect 217318 162596 217324 162648
rect 217376 162636 217382 162648
rect 258166 162636 258172 162648
rect 217376 162608 258172 162636
rect 217376 162596 217382 162608
rect 258166 162596 258172 162608
rect 258224 162596 258230 162648
rect 376294 162596 376300 162648
rect 376352 162636 376358 162648
rect 418706 162636 418712 162648
rect 376352 162608 418712 162636
rect 376352 162596 376358 162608
rect 418706 162596 418712 162608
rect 418764 162596 418770 162648
rect 376478 162528 376484 162580
rect 376536 162568 376542 162580
rect 379238 162568 379244 162580
rect 376536 162540 379244 162568
rect 376536 162528 376542 162540
rect 379238 162528 379244 162540
rect 379296 162568 379302 162580
rect 419534 162568 419540 162580
rect 379296 162540 419540 162568
rect 379296 162528 379302 162540
rect 419534 162528 419540 162540
rect 419592 162528 419598 162580
rect 376570 162460 376576 162512
rect 376628 162500 376634 162512
rect 379790 162500 379796 162512
rect 376628 162472 379796 162500
rect 376628 162460 376634 162472
rect 379790 162460 379796 162472
rect 379848 162460 379854 162512
rect 214650 162392 214656 162444
rect 214708 162432 214714 162444
rect 215754 162432 215760 162444
rect 214708 162404 215760 162432
rect 214708 162392 214714 162404
rect 215754 162392 215760 162404
rect 215812 162432 215818 162444
rect 219342 162432 219348 162444
rect 215812 162404 219348 162432
rect 215812 162392 215818 162404
rect 219342 162392 219348 162404
rect 219400 162392 219406 162444
rect 379606 162256 379612 162308
rect 379664 162296 379670 162308
rect 418154 162296 418160 162308
rect 379664 162268 418160 162296
rect 379664 162256 379670 162268
rect 418154 162256 418160 162268
rect 418212 162256 418218 162308
rect 52086 162188 52092 162240
rect 52144 162228 52150 162240
rect 112070 162228 112076 162240
rect 52144 162200 112076 162228
rect 52144 162188 52150 162200
rect 112070 162188 112076 162200
rect 112128 162188 112134 162240
rect 373534 162188 373540 162240
rect 373592 162228 373598 162240
rect 376202 162228 376208 162240
rect 373592 162200 376208 162228
rect 373592 162188 373598 162200
rect 376202 162188 376208 162200
rect 376260 162228 376266 162240
rect 420914 162228 420920 162240
rect 376260 162200 420920 162228
rect 376260 162188 376266 162200
rect 420914 162188 420920 162200
rect 420972 162188 420978 162240
rect 50890 162120 50896 162172
rect 50948 162160 50954 162172
rect 115750 162160 115756 162172
rect 50948 162132 115756 162160
rect 50948 162120 50954 162132
rect 115750 162120 115756 162132
rect 115808 162120 115814 162172
rect 266354 162160 266360 162172
rect 219406 162132 266360 162160
rect 219158 161780 219164 161832
rect 219216 161820 219222 161832
rect 219406 161820 219434 162132
rect 266354 162120 266360 162132
rect 266412 162120 266418 162172
rect 372338 162120 372344 162172
rect 372396 162160 372402 162172
rect 375006 162160 375012 162172
rect 372396 162132 375012 162160
rect 372396 162120 372402 162132
rect 375006 162120 375012 162132
rect 375064 162160 375070 162172
rect 430574 162160 430580 162172
rect 375064 162132 430580 162160
rect 375064 162120 375070 162132
rect 430574 162120 430580 162132
rect 430632 162120 430638 162172
rect 219526 161820 219532 161832
rect 219216 161792 219532 161820
rect 219216 161780 219222 161792
rect 219526 161780 219532 161792
rect 219584 161780 219590 161832
rect 218974 161508 218980 161560
rect 219032 161548 219038 161560
rect 236638 161548 236644 161560
rect 219032 161520 236644 161548
rect 219032 161508 219038 161520
rect 236638 161508 236644 161520
rect 236696 161508 236702 161560
rect 217870 161440 217876 161492
rect 217928 161480 217934 161492
rect 235258 161480 235264 161492
rect 217928 161452 218468 161480
rect 217928 161440 217934 161452
rect 218440 161412 218468 161452
rect 219084 161452 235264 161480
rect 219084 161412 219112 161452
rect 235258 161440 235264 161452
rect 235316 161440 235322 161492
rect 378962 161440 378968 161492
rect 379020 161480 379026 161492
rect 396718 161480 396724 161492
rect 379020 161452 396724 161480
rect 379020 161440 379026 161452
rect 396718 161440 396724 161452
rect 396776 161440 396782 161492
rect 218440 161384 219112 161412
rect 58710 148996 58716 149048
rect 58768 149036 58774 149048
rect 106274 149036 106280 149048
rect 58768 149008 106280 149036
rect 58768 148996 58774 149008
rect 106274 148996 106280 149008
rect 106332 148996 106338 149048
rect 213546 148996 213552 149048
rect 213604 149036 213610 149048
rect 274726 149036 274732 149048
rect 213604 149008 274732 149036
rect 213604 148996 213610 149008
rect 274726 148996 274732 149008
rect 274784 148996 274790 149048
rect 373810 148996 373816 149048
rect 373868 149036 373874 149048
rect 401594 149036 401600 149048
rect 373868 149008 401600 149036
rect 373868 148996 373874 149008
rect 401594 148996 401600 149008
rect 401652 148996 401658 149048
rect 216306 148928 216312 148980
rect 216364 148968 216370 148980
rect 277394 148968 277400 148980
rect 216364 148940 277400 148968
rect 216364 148928 216370 148940
rect 277394 148928 277400 148940
rect 277452 148928 277458 148980
rect 371602 148928 371608 148980
rect 371660 148968 371666 148980
rect 372430 148968 372436 148980
rect 371660 148940 372436 148968
rect 371660 148928 371666 148940
rect 372430 148928 372436 148940
rect 372488 148968 372494 148980
rect 400214 148968 400220 148980
rect 372488 148940 400220 148968
rect 372488 148928 372494 148940
rect 400214 148928 400220 148940
rect 400272 148928 400278 148980
rect 46566 148792 46572 148844
rect 46624 148832 46630 148844
rect 54938 148832 54944 148844
rect 46624 148804 54944 148832
rect 46624 148792 46630 148804
rect 54938 148792 54944 148804
rect 54996 148832 55002 148844
rect 80054 148832 80060 148844
rect 54996 148804 80060 148832
rect 54996 148792 55002 148804
rect 80054 148792 80060 148804
rect 80112 148792 80118 148844
rect 47854 148724 47860 148776
rect 47912 148764 47918 148776
rect 53466 148764 53472 148776
rect 47912 148736 53472 148764
rect 47912 148724 47918 148736
rect 53466 148724 53472 148736
rect 53524 148764 53530 148776
rect 78674 148764 78680 148776
rect 53524 148736 78680 148764
rect 53524 148724 53530 148736
rect 78674 148724 78680 148736
rect 78732 148724 78738 148776
rect 49050 148656 49056 148708
rect 49108 148696 49114 148708
rect 51994 148696 52000 148708
rect 49108 148668 52000 148696
rect 49108 148656 49114 148668
rect 51994 148656 52000 148668
rect 52052 148696 52058 148708
rect 81434 148696 81440 148708
rect 52052 148668 81440 148696
rect 52052 148656 52058 148668
rect 81434 148656 81440 148668
rect 81492 148656 81498 148708
rect 52914 148588 52920 148640
rect 52972 148628 52978 148640
rect 55858 148628 55864 148640
rect 52972 148600 55864 148628
rect 52972 148588 52978 148600
rect 55858 148588 55864 148600
rect 55916 148628 55922 148640
rect 100018 148628 100024 148640
rect 55916 148600 100024 148628
rect 55916 148588 55922 148600
rect 100018 148588 100024 148600
rect 100076 148588 100082 148640
rect 213270 148588 213276 148640
rect 213328 148628 213334 148640
rect 238754 148628 238760 148640
rect 213328 148600 238760 148628
rect 213328 148588 213334 148600
rect 238754 148588 238760 148600
rect 238812 148588 238818 148640
rect 46106 148520 46112 148572
rect 46164 148560 46170 148572
rect 59814 148560 59820 148572
rect 46164 148532 59820 148560
rect 46164 148520 46170 148532
rect 59814 148520 59820 148532
rect 59872 148560 59878 148572
rect 107654 148560 107660 148572
rect 59872 148532 107660 148560
rect 59872 148520 59878 148532
rect 107654 148520 107660 148532
rect 107712 148520 107718 148572
rect 214926 148520 214932 148572
rect 214984 148560 214990 148572
rect 240134 148560 240140 148572
rect 214984 148532 240140 148560
rect 214984 148520 214990 148532
rect 240134 148520 240140 148532
rect 240192 148520 240198 148572
rect 59170 148452 59176 148504
rect 59228 148492 59234 148504
rect 107746 148492 107752 148504
rect 59228 148464 107752 148492
rect 59228 148452 59234 148464
rect 107746 148452 107752 148464
rect 107804 148452 107810 148504
rect 213730 148452 213736 148504
rect 213788 148492 213794 148504
rect 241514 148492 241520 148504
rect 213788 148464 241520 148492
rect 213788 148452 213794 148464
rect 241514 148452 241520 148464
rect 241572 148452 241578 148504
rect 374730 148452 374736 148504
rect 374788 148492 374794 148504
rect 397454 148492 397460 148504
rect 374788 148464 397460 148492
rect 374788 148452 374794 148464
rect 397454 148452 397460 148464
rect 397512 148452 397518 148504
rect 53558 148384 53564 148436
rect 53616 148424 53622 148436
rect 114646 148424 114652 148436
rect 53616 148396 114652 148424
rect 53616 148384 53622 148396
rect 114646 148384 114652 148396
rect 114704 148384 114710 148436
rect 213086 148384 213092 148436
rect 213144 148424 213150 148436
rect 215018 148424 215024 148436
rect 213144 148396 215024 148424
rect 213144 148384 213150 148396
rect 215018 148384 215024 148396
rect 215076 148424 215082 148436
rect 270494 148424 270500 148436
rect 215076 148396 270500 148424
rect 215076 148384 215082 148396
rect 270494 148384 270500 148396
rect 270552 148384 270558 148436
rect 374822 148384 374828 148436
rect 374880 148424 374886 148436
rect 398834 148424 398840 148436
rect 374880 148396 398840 148424
rect 374880 148384 374886 148396
rect 398834 148384 398840 148396
rect 398892 148384 398898 148436
rect 53098 148316 53104 148368
rect 53156 148356 53162 148368
rect 114738 148356 114744 148368
rect 53156 148328 114744 148356
rect 53156 148316 53162 148328
rect 114738 148316 114744 148328
rect 114796 148316 114802 148368
rect 213454 148316 213460 148368
rect 213512 148356 213518 148368
rect 215938 148356 215944 148368
rect 213512 148328 215944 148356
rect 213512 148316 213518 148328
rect 215938 148316 215944 148328
rect 215996 148356 216002 148368
rect 271874 148356 271880 148368
rect 215996 148328 271880 148356
rect 215996 148316 216002 148328
rect 271874 148316 271880 148328
rect 271932 148316 271938 148368
rect 373074 148316 373080 148368
rect 373132 148356 373138 148368
rect 375190 148356 375196 148368
rect 373132 148328 375196 148356
rect 373132 148316 373138 148328
rect 375190 148316 375196 148328
rect 375248 148356 375254 148368
rect 434714 148356 434720 148368
rect 375248 148328 434720 148356
rect 375248 148316 375254 148328
rect 434714 148316 434720 148328
rect 434772 148316 434778 148368
rect 48222 147568 48228 147620
rect 48280 147608 48286 147620
rect 58894 147608 58900 147620
rect 48280 147580 58900 147608
rect 48280 147568 48286 147580
rect 58894 147568 58900 147580
rect 58952 147608 58958 147620
rect 59170 147608 59176 147620
rect 58952 147580 59176 147608
rect 58952 147568 58958 147580
rect 59170 147568 59176 147580
rect 59228 147568 59234 147620
rect 210878 147568 210884 147620
rect 210936 147608 210942 147620
rect 214558 147608 214564 147620
rect 210936 147580 214564 147608
rect 210936 147568 210942 147580
rect 214558 147568 214564 147580
rect 214616 147608 214622 147620
rect 214926 147608 214932 147620
rect 214616 147580 214932 147608
rect 214616 147568 214622 147580
rect 214926 147568 214932 147580
rect 214984 147568 214990 147620
rect 371050 147568 371056 147620
rect 371108 147608 371114 147620
rect 374730 147608 374736 147620
rect 371108 147580 374736 147608
rect 371108 147568 371114 147580
rect 374730 147568 374736 147580
rect 374788 147568 374794 147620
rect 212350 147500 212356 147552
rect 212408 147540 212414 147552
rect 213270 147540 213276 147552
rect 212408 147512 213276 147540
rect 212408 147500 212414 147512
rect 213270 147500 213276 147512
rect 213328 147500 213334 147552
rect 368290 147500 368296 147552
rect 368348 147540 368354 147552
rect 374822 147540 374828 147552
rect 368348 147512 374828 147540
rect 368348 147500 368354 147512
rect 374822 147500 374828 147512
rect 374880 147500 374886 147552
rect 208302 147432 208308 147484
rect 208360 147472 208366 147484
rect 213178 147472 213184 147484
rect 208360 147444 213184 147472
rect 208360 147432 208366 147444
rect 213178 147432 213184 147444
rect 213236 147472 213242 147484
rect 213730 147472 213736 147484
rect 213236 147444 213736 147472
rect 213236 147432 213242 147444
rect 213730 147432 213736 147444
rect 213788 147432 213794 147484
rect 59004 146288 59492 146316
rect 48038 146208 48044 146260
rect 48096 146248 48102 146260
rect 51718 146248 51724 146260
rect 48096 146220 51724 146248
rect 48096 146208 48102 146220
rect 51718 146208 51724 146220
rect 51776 146208 51782 146260
rect 56962 146208 56968 146260
rect 57020 146248 57026 146260
rect 57238 146248 57244 146260
rect 57020 146220 57244 146248
rect 57020 146208 57026 146220
rect 57238 146208 57244 146220
rect 57296 146248 57302 146260
rect 59004 146248 59032 146288
rect 57296 146220 59032 146248
rect 57296 146208 57302 146220
rect 59078 146208 59084 146260
rect 59136 146248 59142 146260
rect 59354 146248 59360 146260
rect 59136 146220 59360 146248
rect 59136 146208 59142 146220
rect 59354 146208 59360 146220
rect 59412 146208 59418 146260
rect 59464 146248 59492 146288
rect 213730 146276 213736 146328
rect 213788 146316 213794 146328
rect 213788 146288 274680 146316
rect 213788 146276 213794 146288
rect 91094 146248 91100 146260
rect 59464 146220 91100 146248
rect 91094 146208 91100 146220
rect 91152 146208 91158 146260
rect 179046 146208 179052 146260
rect 179104 146248 179110 146260
rect 197630 146248 197636 146260
rect 179104 146220 197636 146248
rect 179104 146208 179110 146220
rect 197630 146208 197636 146220
rect 197688 146208 197694 146260
rect 235994 146248 236000 146260
rect 219406 146220 236000 146248
rect 53190 146140 53196 146192
rect 53248 146180 53254 146192
rect 86954 146180 86960 146192
rect 53248 146152 86960 146180
rect 53248 146140 53254 146152
rect 86954 146140 86960 146152
rect 87012 146140 87018 146192
rect 179690 146140 179696 146192
rect 179748 146180 179754 146192
rect 197538 146180 197544 146192
rect 179748 146152 197544 146180
rect 179748 146140 179754 146152
rect 197538 146140 197544 146152
rect 197596 146140 197602 146192
rect 214466 146140 214472 146192
rect 214524 146180 214530 146192
rect 215846 146180 215852 146192
rect 214524 146152 215852 146180
rect 214524 146140 214530 146152
rect 215846 146140 215852 146152
rect 215904 146180 215910 146192
rect 219406 146180 219434 146220
rect 235994 146208 236000 146220
rect 236052 146208 236058 146260
rect 236638 146208 236644 146260
rect 236696 146248 236702 146260
rect 256694 146248 256700 146260
rect 236696 146220 256700 146248
rect 236696 146208 236702 146220
rect 256694 146208 256700 146220
rect 256752 146208 256758 146260
rect 274652 146248 274680 146288
rect 274818 146248 274824 146260
rect 274652 146220 274824 146248
rect 274818 146208 274824 146220
rect 274876 146248 274882 146260
rect 356790 146248 356796 146260
rect 274876 146220 356796 146248
rect 274876 146208 274882 146220
rect 356790 146208 356796 146220
rect 356848 146208 356854 146260
rect 377582 146208 377588 146260
rect 377640 146248 377646 146260
rect 378042 146248 378048 146260
rect 377640 146220 378048 146248
rect 377640 146208 377646 146220
rect 378042 146208 378048 146220
rect 378100 146208 378106 146260
rect 378594 146208 378600 146260
rect 378652 146248 378658 146260
rect 379330 146248 379336 146260
rect 378652 146220 379336 146248
rect 378652 146208 378658 146220
rect 379330 146208 379336 146220
rect 379388 146208 379394 146260
rect 403066 146248 403072 146260
rect 383626 146220 403072 146248
rect 215904 146152 219434 146180
rect 215904 146140 215910 146152
rect 235258 146140 235264 146192
rect 235316 146180 235322 146192
rect 255406 146180 255412 146192
rect 235316 146152 255412 146180
rect 235316 146140 235322 146152
rect 255406 146140 255412 146152
rect 255464 146140 255470 146192
rect 338482 146140 338488 146192
rect 338540 146180 338546 146192
rect 360194 146180 360200 146192
rect 338540 146152 360200 146180
rect 338540 146140 338546 146152
rect 360194 146140 360200 146152
rect 360252 146140 360258 146192
rect 377398 146140 377404 146192
rect 377456 146180 377462 146192
rect 377950 146180 377956 146192
rect 377456 146152 377956 146180
rect 377456 146140 377462 146152
rect 377950 146140 377956 146152
rect 378008 146140 378014 146192
rect 383626 146180 383654 146220
rect 403066 146208 403072 146220
rect 403124 146208 403130 146260
rect 379164 146152 383654 146180
rect 58618 146072 58624 146124
rect 58676 146112 58682 146124
rect 59170 146112 59176 146124
rect 58676 146084 59176 146112
rect 58676 146072 58682 146084
rect 59170 146072 59176 146084
rect 59228 146072 59234 146124
rect 59722 146072 59728 146124
rect 59780 146112 59786 146124
rect 60734 146112 60740 146124
rect 59780 146084 60740 146112
rect 59780 146072 59786 146084
rect 60734 146072 60740 146084
rect 60792 146112 60798 146124
rect 66254 146112 66260 146124
rect 60792 146084 66260 146112
rect 60792 146072 60798 146084
rect 66254 146072 66260 146084
rect 66312 146072 66318 146124
rect 92474 146112 92480 146124
rect 66364 146084 92480 146112
rect 59354 146004 59360 146056
rect 59412 146044 59418 146056
rect 66364 146044 66392 146084
rect 92474 146072 92480 146084
rect 92532 146072 92538 146124
rect 219250 146072 219256 146124
rect 219308 146112 219314 146124
rect 251174 146112 251180 146124
rect 219308 146084 251180 146112
rect 219308 146072 219314 146084
rect 251174 146072 251180 146084
rect 251232 146072 251238 146124
rect 340230 146072 340236 146124
rect 340288 146112 340294 146124
rect 357618 146112 357624 146124
rect 340288 146084 357624 146112
rect 340288 146072 340294 146084
rect 357618 146072 357624 146084
rect 357676 146072 357682 146124
rect 375926 146072 375932 146124
rect 375984 146112 375990 146124
rect 378502 146112 378508 146124
rect 375984 146084 378508 146112
rect 375984 146072 375990 146084
rect 378502 146072 378508 146084
rect 378560 146112 378566 146124
rect 379164 146112 379192 146152
rect 396718 146140 396724 146192
rect 396776 146180 396782 146192
rect 416774 146180 416780 146192
rect 396776 146152 416780 146180
rect 396776 146140 396782 146152
rect 416774 146140 416780 146152
rect 416832 146140 416838 146192
rect 500218 146140 500224 146192
rect 500276 146180 500282 146192
rect 517514 146180 517520 146192
rect 500276 146152 517520 146180
rect 500276 146140 500282 146152
rect 517514 146140 517520 146152
rect 517572 146180 517578 146192
rect 517698 146180 517704 146192
rect 517572 146152 517704 146180
rect 517572 146140 517578 146152
rect 517698 146140 517704 146152
rect 517756 146140 517762 146192
rect 378560 146084 379192 146112
rect 378560 146072 378566 146084
rect 379238 146072 379244 146124
rect 379296 146112 379302 146124
rect 379974 146112 379980 146124
rect 379296 146084 379980 146112
rect 379296 146072 379302 146084
rect 379974 146072 379980 146084
rect 380032 146112 380038 146124
rect 412634 146112 412640 146124
rect 380032 146084 412640 146112
rect 380032 146072 380038 146084
rect 412634 146072 412640 146084
rect 412692 146072 412698 146124
rect 498654 146072 498660 146124
rect 498712 146112 498718 146124
rect 517790 146112 517796 146124
rect 498712 146084 517796 146112
rect 498712 146072 498718 146084
rect 517790 146072 517796 146084
rect 517848 146072 517854 146124
rect 59412 146016 66392 146044
rect 59412 146004 59418 146016
rect 66438 146004 66444 146056
rect 66496 146044 66502 146056
rect 93854 146044 93860 146056
rect 66496 146016 93860 146044
rect 66496 146004 66502 146016
rect 93854 146004 93860 146016
rect 93912 146004 93918 146056
rect 215754 146004 215760 146056
rect 215812 146044 215818 146056
rect 217962 146044 217968 146056
rect 215812 146016 217968 146044
rect 215812 146004 215818 146016
rect 217962 146004 217968 146016
rect 218020 146044 218026 146056
rect 249886 146044 249892 146056
rect 218020 146016 249892 146044
rect 218020 146004 218026 146016
rect 249886 146004 249892 146016
rect 249944 146004 249950 146056
rect 379330 146004 379336 146056
rect 379388 146044 379394 146056
rect 411254 146044 411260 146056
rect 379388 146016 411260 146044
rect 379388 146004 379394 146016
rect 411254 146004 411260 146016
rect 411312 146004 411318 146056
rect 56134 145936 56140 145988
rect 56192 145976 56198 145988
rect 88426 145976 88432 145988
rect 56192 145948 88432 145976
rect 56192 145936 56198 145948
rect 88426 145936 88432 145948
rect 88484 145936 88490 145988
rect 218422 145936 218428 145988
rect 218480 145976 218486 145988
rect 219802 145976 219808 145988
rect 218480 145948 219808 145976
rect 218480 145936 218486 145948
rect 219802 145936 219808 145948
rect 219860 145936 219866 145988
rect 219894 145936 219900 145988
rect 219952 145936 219958 145988
rect 251266 145976 251272 145988
rect 221936 145948 251272 145976
rect 59170 145868 59176 145920
rect 59228 145908 59234 145920
rect 89806 145908 89812 145920
rect 59228 145880 89812 145908
rect 59228 145868 59234 145880
rect 89806 145868 89812 145880
rect 89864 145868 89870 145920
rect 217042 145868 217048 145920
rect 217100 145908 217106 145920
rect 219912 145908 219940 145936
rect 221936 145908 221964 145948
rect 251266 145936 251272 145948
rect 251324 145936 251330 145988
rect 377950 145936 377956 145988
rect 378008 145936 378014 145988
rect 378042 145936 378048 145988
rect 378100 145976 378106 145988
rect 379146 145976 379152 145988
rect 378100 145948 379152 145976
rect 378100 145936 378106 145948
rect 379146 145936 379152 145948
rect 379204 145976 379210 145988
rect 409966 145976 409972 145988
rect 379204 145948 409972 145976
rect 379204 145936 379210 145948
rect 409966 145936 409972 145948
rect 410024 145936 410030 145988
rect 217100 145880 221964 145908
rect 217100 145868 217106 145880
rect 224218 145868 224224 145920
rect 224276 145908 224282 145920
rect 244274 145908 244280 145920
rect 224276 145880 244280 145908
rect 224276 145868 224282 145880
rect 244274 145868 244280 145880
rect 244332 145868 244338 145920
rect 374546 145868 374552 145920
rect 374604 145908 374610 145920
rect 374822 145908 374828 145920
rect 374604 145880 374828 145908
rect 374604 145868 374610 145880
rect 374822 145868 374828 145880
rect 374880 145868 374886 145920
rect 377968 145908 377996 145936
rect 408494 145908 408500 145920
rect 377968 145880 408500 145908
rect 408494 145868 408500 145880
rect 408552 145868 408558 145920
rect 54570 145800 54576 145852
rect 54628 145840 54634 145852
rect 54846 145840 54852 145852
rect 54628 145812 54852 145840
rect 54628 145800 54634 145812
rect 54846 145800 54852 145812
rect 54904 145840 54910 145852
rect 85574 145840 85580 145852
rect 54904 145812 85580 145840
rect 54904 145800 54910 145812
rect 85574 145800 85580 145812
rect 85632 145800 85638 145852
rect 216122 145800 216128 145852
rect 216180 145840 216186 145852
rect 216858 145840 216864 145852
rect 216180 145812 216864 145840
rect 216180 145800 216186 145812
rect 216858 145800 216864 145812
rect 216916 145840 216922 145852
rect 247126 145840 247132 145852
rect 216916 145812 247132 145840
rect 216916 145800 216922 145812
rect 247126 145800 247132 145812
rect 247184 145800 247190 145852
rect 374840 145840 374868 145868
rect 404354 145840 404360 145852
rect 374840 145812 404360 145840
rect 404354 145800 404360 145812
rect 404412 145800 404418 145852
rect 58710 145732 58716 145784
rect 58768 145772 58774 145784
rect 84194 145772 84200 145784
rect 58768 145744 84200 145772
rect 58768 145732 58774 145744
rect 84194 145732 84200 145744
rect 84252 145732 84258 145784
rect 218146 145732 218152 145784
rect 218204 145772 218210 145784
rect 218882 145772 218888 145784
rect 218204 145744 218888 145772
rect 218204 145732 218210 145744
rect 218882 145732 218888 145744
rect 218940 145772 218946 145784
rect 245654 145772 245660 145784
rect 218940 145744 245660 145772
rect 218940 145732 218946 145744
rect 245654 145732 245660 145744
rect 245712 145732 245718 145784
rect 374546 145732 374552 145784
rect 374604 145772 374610 145784
rect 375650 145772 375656 145784
rect 374604 145744 375656 145772
rect 374604 145732 374610 145744
rect 375650 145732 375656 145744
rect 375708 145772 375714 145784
rect 402974 145772 402980 145784
rect 375708 145744 402980 145772
rect 375708 145732 375714 145744
rect 402974 145732 402980 145744
rect 403032 145732 403038 145784
rect 56410 145664 56416 145716
rect 56468 145704 56474 145716
rect 84286 145704 84292 145716
rect 56468 145676 84292 145704
rect 56468 145664 56474 145676
rect 84286 145664 84292 145676
rect 84344 145664 84350 145716
rect 216214 145664 216220 145716
rect 216272 145704 216278 145716
rect 216490 145704 216496 145716
rect 216272 145676 216496 145704
rect 216272 145664 216278 145676
rect 216490 145664 216496 145676
rect 216548 145704 216554 145716
rect 242894 145704 242900 145716
rect 216548 145676 242900 145704
rect 216548 145664 216554 145676
rect 242894 145664 242900 145676
rect 242952 145664 242958 145716
rect 378778 145664 378784 145716
rect 378836 145704 378842 145716
rect 407206 145704 407212 145716
rect 378836 145676 407212 145704
rect 378836 145664 378842 145676
rect 407206 145664 407212 145676
rect 407264 145664 407270 145716
rect 50062 145596 50068 145648
rect 50120 145636 50126 145648
rect 54386 145636 54392 145648
rect 50120 145608 54392 145636
rect 50120 145596 50126 145608
rect 54386 145596 54392 145608
rect 54444 145636 54450 145648
rect 82814 145636 82820 145648
rect 54444 145608 82820 145636
rect 54444 145596 54450 145608
rect 82814 145596 82820 145608
rect 82872 145596 82878 145648
rect 214834 145596 214840 145648
rect 214892 145636 214898 145648
rect 224218 145636 224224 145648
rect 214892 145608 224224 145636
rect 214892 145596 214898 145608
rect 224218 145596 224224 145608
rect 224276 145596 224282 145648
rect 224310 145596 224316 145648
rect 224368 145636 224374 145648
rect 244366 145636 244372 145648
rect 224368 145608 244372 145636
rect 224368 145596 224374 145608
rect 244366 145596 244372 145608
rect 244424 145596 244430 145648
rect 376386 145596 376392 145648
rect 376444 145636 376450 145648
rect 405734 145636 405740 145648
rect 376444 145608 405740 145636
rect 376444 145596 376450 145608
rect 405734 145596 405740 145608
rect 405792 145596 405798 145648
rect 517514 145596 517520 145648
rect 517572 145636 517578 145648
rect 580258 145636 580264 145648
rect 517572 145608 580264 145636
rect 517572 145596 517578 145608
rect 580258 145596 580264 145608
rect 580316 145596 580322 145648
rect 58618 145528 58624 145580
rect 58676 145568 58682 145580
rect 91186 145568 91192 145580
rect 58676 145540 91192 145568
rect 58676 145528 58682 145540
rect 91186 145528 91192 145540
rect 91244 145528 91250 145580
rect 191282 145528 191288 145580
rect 191340 145568 191346 145580
rect 201494 145568 201500 145580
rect 191340 145540 201500 145568
rect 191340 145528 191346 145540
rect 201494 145528 201500 145540
rect 201552 145568 201558 145580
rect 204898 145568 204904 145580
rect 201552 145540 204904 145568
rect 201552 145528 201558 145540
rect 204898 145528 204904 145540
rect 204956 145528 204962 145580
rect 216950 145528 216956 145580
rect 217008 145568 217014 145580
rect 248414 145568 248420 145580
rect 217008 145540 248420 145568
rect 217008 145528 217014 145540
rect 248414 145528 248420 145540
rect 248472 145528 248478 145580
rect 280062 145528 280068 145580
rect 280120 145568 280126 145580
rect 307662 145568 307668 145580
rect 280120 145540 307668 145568
rect 280120 145528 280126 145540
rect 307662 145528 307668 145540
rect 307720 145528 307726 145580
rect 351638 145528 351644 145580
rect 351696 145568 351702 145580
rect 358078 145568 358084 145580
rect 351696 145540 358084 145568
rect 351696 145528 351702 145540
rect 358078 145528 358084 145540
rect 358136 145568 358142 145580
rect 358722 145568 358728 145580
rect 358136 145540 358728 145568
rect 358136 145528 358142 145540
rect 358722 145528 358728 145540
rect 358780 145568 358786 145580
rect 510522 145568 510528 145580
rect 358780 145540 510528 145568
rect 358780 145528 358786 145540
rect 510522 145528 510528 145540
rect 510580 145528 510586 145580
rect 517790 145528 517796 145580
rect 517848 145568 517854 145580
rect 580350 145568 580356 145580
rect 517848 145540 580356 145568
rect 517848 145528 517854 145540
rect 580350 145528 580356 145540
rect 580408 145528 580414 145580
rect 51718 145460 51724 145512
rect 51776 145500 51782 145512
rect 77294 145500 77300 145512
rect 51776 145472 77300 145500
rect 51776 145460 51782 145472
rect 77294 145460 77300 145472
rect 77352 145460 77358 145512
rect 218514 145460 218520 145512
rect 218572 145500 218578 145512
rect 236086 145500 236092 145512
rect 218572 145472 236092 145500
rect 218572 145460 218578 145472
rect 236086 145460 236092 145472
rect 236144 145460 236150 145512
rect 378686 145460 378692 145512
rect 378744 145500 378750 145512
rect 396074 145500 396080 145512
rect 378744 145472 396080 145500
rect 378744 145460 378750 145472
rect 396074 145460 396080 145472
rect 396132 145460 396138 145512
rect 48130 145392 48136 145444
rect 48188 145432 48194 145444
rect 54478 145432 54484 145444
rect 48188 145404 54484 145432
rect 48188 145392 48194 145404
rect 54478 145392 54484 145404
rect 54536 145432 54542 145444
rect 75914 145432 75920 145444
rect 54536 145404 75920 145432
rect 54536 145392 54542 145404
rect 75914 145392 75920 145404
rect 75972 145392 75978 145444
rect 219710 145392 219716 145444
rect 219768 145432 219774 145444
rect 253934 145432 253940 145444
rect 219768 145404 253940 145432
rect 219768 145392 219774 145404
rect 253934 145392 253940 145404
rect 253992 145392 253998 145444
rect 378870 145392 378876 145444
rect 378928 145432 378934 145444
rect 396166 145432 396172 145444
rect 378928 145404 396172 145432
rect 378928 145392 378934 145404
rect 396166 145392 396172 145404
rect 396224 145392 396230 145444
rect 46658 145324 46664 145376
rect 46716 145364 46722 145376
rect 54754 145364 54760 145376
rect 46716 145336 54760 145364
rect 46716 145324 46722 145336
rect 54754 145324 54760 145336
rect 54812 145364 54818 145376
rect 76006 145364 76012 145376
rect 54812 145336 76012 145364
rect 54812 145324 54818 145336
rect 76006 145324 76012 145336
rect 76064 145324 76070 145376
rect 219802 145324 219808 145376
rect 219860 145364 219866 145376
rect 252646 145364 252652 145376
rect 219860 145336 252652 145364
rect 219860 145324 219866 145336
rect 252646 145324 252652 145336
rect 252704 145324 252710 145376
rect 379882 145324 379888 145376
rect 379940 145364 379946 145376
rect 414014 145364 414020 145376
rect 379940 145336 414020 145364
rect 379940 145324 379946 145336
rect 414014 145324 414020 145336
rect 414072 145324 414078 145376
rect 377582 145256 377588 145308
rect 377640 145296 377646 145308
rect 411346 145296 411352 145308
rect 377640 145268 411352 145296
rect 377640 145256 377646 145268
rect 411346 145256 411352 145268
rect 411404 145256 411410 145308
rect 216030 144984 216036 145036
rect 216088 145024 216094 145036
rect 224310 145024 224316 145036
rect 216088 144996 224316 145024
rect 216088 144984 216094 144996
rect 224310 144984 224316 144996
rect 224368 144984 224374 145036
rect 377398 144956 377404 144968
rect 376496 144928 377404 144956
rect 54662 144848 54668 144900
rect 54720 144888 54726 144900
rect 56042 144888 56048 144900
rect 54720 144860 56048 144888
rect 54720 144848 54726 144860
rect 56042 144848 56048 144860
rect 56100 144888 56106 144900
rect 56410 144888 56416 144900
rect 56100 144860 56416 144888
rect 56100 144848 56106 144860
rect 56410 144848 56416 144860
rect 56468 144848 56474 144900
rect 214282 144848 214288 144900
rect 214340 144888 214346 144900
rect 216950 144888 216956 144900
rect 214340 144860 216956 144888
rect 214340 144848 214346 144860
rect 216950 144848 216956 144860
rect 217008 144888 217014 144900
rect 217134 144888 217140 144900
rect 217008 144860 217140 144888
rect 217008 144848 217014 144860
rect 217134 144848 217140 144860
rect 217192 144848 217198 144900
rect 307662 144848 307668 144900
rect 307720 144888 307726 144900
rect 356606 144888 356612 144900
rect 307720 144860 356612 144888
rect 307720 144848 307726 144860
rect 356606 144848 356612 144860
rect 356664 144848 356670 144900
rect 51810 144780 51816 144832
rect 51868 144820 51874 144832
rect 58710 144820 58716 144832
rect 51868 144792 58716 144820
rect 51868 144780 51874 144792
rect 58710 144780 58716 144792
rect 58768 144780 58774 144832
rect 209406 144780 209412 144832
rect 209464 144820 209470 144832
rect 213454 144820 213460 144832
rect 209464 144792 213460 144820
rect 209464 144780 209470 144792
rect 213454 144780 213460 144792
rect 213512 144780 213518 144832
rect 373902 144780 373908 144832
rect 373960 144820 373966 144832
rect 376018 144820 376024 144832
rect 373960 144792 376024 144820
rect 373960 144780 373966 144792
rect 376018 144780 376024 144792
rect 376076 144820 376082 144832
rect 376386 144820 376392 144832
rect 376076 144792 376392 144820
rect 376076 144780 376082 144792
rect 376386 144780 376392 144792
rect 376444 144780 376450 144832
rect 53282 144712 53288 144764
rect 53340 144752 53346 144764
rect 58618 144752 58624 144764
rect 53340 144724 58624 144752
rect 53340 144712 53346 144724
rect 58618 144712 58624 144724
rect 58676 144712 58682 144764
rect 212994 144712 213000 144764
rect 213052 144752 213058 144764
rect 216030 144752 216036 144764
rect 213052 144724 216036 144752
rect 213052 144712 213058 144724
rect 216030 144712 216036 144724
rect 216088 144712 216094 144764
rect 376496 144752 376524 144928
rect 377398 144916 377404 144928
rect 377456 144916 377462 144968
rect 376404 144724 376524 144752
rect 376404 144696 376432 144724
rect 47578 144644 47584 144696
rect 47636 144684 47642 144696
rect 55950 144684 55956 144696
rect 47636 144656 55956 144684
rect 47636 144644 47642 144656
rect 55950 144644 55956 144656
rect 56008 144684 56014 144696
rect 56318 144684 56324 144696
rect 56008 144656 56324 144684
rect 56008 144644 56014 144656
rect 56318 144644 56324 144656
rect 56376 144644 56382 144696
rect 376386 144644 376392 144696
rect 376444 144644 376450 144696
rect 56226 144576 56232 144628
rect 56284 144616 56290 144628
rect 56284 144588 56364 144616
rect 56284 144576 56290 144588
rect 56336 144424 56364 144588
rect 375742 144576 375748 144628
rect 375800 144616 375806 144628
rect 378778 144616 378784 144628
rect 375800 144588 378784 144616
rect 375800 144576 375806 144588
rect 378778 144576 378784 144588
rect 378836 144576 378842 144628
rect 56318 144372 56324 144424
rect 56376 144372 56382 144424
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 21358 97968 21364 97980
rect 3568 97940 21364 97968
rect 3568 97928 3574 97940
rect 21358 97928 21364 97940
rect 21416 97928 21422 97980
rect 520182 79976 520188 80028
rect 520240 80016 520246 80028
rect 580442 80016 580448 80028
rect 520240 79988 580448 80016
rect 520240 79976 520246 79988
rect 580442 79976 580448 79988
rect 580500 79976 580506 80028
rect 42610 70320 42616 70372
rect 42668 70360 42674 70372
rect 57606 70360 57612 70372
rect 42668 70332 57612 70360
rect 42668 70320 42674 70332
rect 57606 70320 57612 70332
rect 57664 70320 57670 70372
rect 209038 70320 209044 70372
rect 209096 70360 209102 70372
rect 216674 70360 216680 70372
rect 209096 70332 216680 70360
rect 209096 70320 209102 70332
rect 216674 70320 216680 70332
rect 216732 70320 216738 70372
rect 362310 70320 362316 70372
rect 362368 70360 362374 70372
rect 376938 70360 376944 70372
rect 362368 70332 376944 70360
rect 362368 70320 362374 70332
rect 376938 70320 376944 70332
rect 376996 70320 377002 70372
rect 358722 68280 358728 68332
rect 358780 68320 358786 68332
rect 376938 68320 376944 68332
rect 358780 68292 376944 68320
rect 358780 68280 358786 68292
rect 376938 68280 376944 68292
rect 376996 68280 377002 68332
rect 358078 68144 358084 68196
rect 358136 68184 358142 68196
rect 358722 68184 358728 68196
rect 358136 68156 358728 68184
rect 358136 68144 358142 68156
rect 358722 68144 358728 68156
rect 358780 68144 358786 68196
rect 204898 67600 204904 67652
rect 204956 67640 204962 67652
rect 216674 67640 216680 67652
rect 204956 67612 216680 67640
rect 204956 67600 204962 67612
rect 216674 67600 216680 67612
rect 216732 67600 216738 67652
rect 54478 59712 54484 59764
rect 54536 59752 54542 59764
rect 77110 59752 77116 59764
rect 54536 59724 77116 59752
rect 54536 59712 54542 59724
rect 77110 59712 77116 59724
rect 77168 59712 77174 59764
rect 378870 59712 378876 59764
rect 378928 59752 378934 59764
rect 397086 59752 397092 59764
rect 378928 59724 397092 59752
rect 378928 59712 378934 59724
rect 397086 59712 397092 59724
rect 397144 59712 397150 59764
rect 54386 59644 54392 59696
rect 54444 59684 54450 59696
rect 83090 59684 83096 59696
rect 54444 59656 83096 59684
rect 54444 59644 54450 59656
rect 83090 59644 83096 59656
rect 83148 59644 83154 59696
rect 218514 59644 218520 59696
rect 218572 59684 218578 59696
rect 235994 59684 236000 59696
rect 218572 59656 236000 59684
rect 218572 59644 218578 59656
rect 235994 59644 236000 59656
rect 236052 59644 236058 59696
rect 378686 59644 378692 59696
rect 378744 59684 378750 59696
rect 396074 59684 396080 59696
rect 378744 59656 396080 59684
rect 378744 59644 378750 59656
rect 396074 59644 396080 59656
rect 396132 59644 396138 59696
rect 58986 59576 58992 59628
rect 59044 59616 59050 59628
rect 100754 59616 100760 59628
rect 59044 59588 100760 59616
rect 59044 59576 59050 59588
rect 100754 59576 100760 59588
rect 100812 59576 100818 59628
rect 214466 59576 214472 59628
rect 214524 59616 214530 59628
rect 237098 59616 237104 59628
rect 214524 59588 237104 59616
rect 214524 59576 214530 59588
rect 237098 59576 237104 59588
rect 237156 59576 237162 59628
rect 374546 59576 374552 59628
rect 374604 59616 374610 59628
rect 403066 59616 403072 59628
rect 374604 59588 403072 59616
rect 374604 59576 374610 59588
rect 403066 59576 403072 59588
rect 403124 59576 403130 59628
rect 54570 59508 54576 59560
rect 54628 59548 54634 59560
rect 101766 59548 101772 59560
rect 54628 59520 101772 59548
rect 54628 59508 54634 59520
rect 101766 59508 101772 59520
rect 101824 59508 101830 59560
rect 217870 59508 217876 59560
rect 217928 59548 217934 59560
rect 255866 59548 255872 59560
rect 217928 59520 255872 59548
rect 217928 59508 217934 59520
rect 255866 59508 255872 59520
rect 255924 59508 255930 59560
rect 378962 59508 378968 59560
rect 379020 59548 379026 59560
rect 416958 59548 416964 59560
rect 379020 59520 416964 59548
rect 379020 59508 379026 59520
rect 416958 59508 416964 59520
rect 417016 59508 417022 59560
rect 58894 59440 58900 59492
rect 58952 59480 58958 59492
rect 107562 59480 107568 59492
rect 58952 59452 107568 59480
rect 58952 59440 58958 59452
rect 107562 59440 107568 59452
rect 107620 59440 107626 59492
rect 218974 59440 218980 59492
rect 219032 59480 219038 59492
rect 256970 59480 256976 59492
rect 219032 59452 256976 59480
rect 219032 59440 219038 59452
rect 256970 59440 256976 59452
rect 257028 59440 257034 59492
rect 377490 59440 377496 59492
rect 377548 59480 377554 59492
rect 423950 59480 423956 59492
rect 377548 59452 423956 59480
rect 377548 59440 377554 59452
rect 423950 59440 423956 59452
rect 424008 59440 424014 59492
rect 52270 59372 52276 59424
rect 52328 59412 52334 59424
rect 113542 59412 113548 59424
rect 52328 59384 113548 59412
rect 52328 59372 52334 59384
rect 113542 59372 113548 59384
rect 113600 59372 113606 59424
rect 216582 59372 216588 59424
rect 216640 59412 216646 59424
rect 262858 59412 262864 59424
rect 216640 59384 262864 59412
rect 216640 59372 216646 59384
rect 262858 59372 262864 59384
rect 262916 59372 262922 59424
rect 376110 59372 376116 59424
rect 376168 59412 376174 59424
rect 422846 59412 422852 59424
rect 376168 59384 422852 59412
rect 376168 59372 376174 59384
rect 422846 59372 422852 59384
rect 422904 59372 422910 59424
rect 56042 59304 56048 59356
rect 56100 59344 56106 59356
rect 84194 59344 84200 59356
rect 56100 59316 84200 59344
rect 56100 59304 56106 59316
rect 84194 59304 84200 59316
rect 84252 59304 84258 59356
rect 217962 59304 217968 59356
rect 218020 59344 218026 59356
rect 358078 59344 358084 59356
rect 218020 59316 358084 59344
rect 218020 59304 218026 59316
rect 358078 59304 358084 59316
rect 358136 59304 358142 59356
rect 379882 59304 379888 59356
rect 379940 59344 379946 59356
rect 414566 59344 414572 59356
rect 379940 59316 414572 59344
rect 379940 59304 379946 59316
rect 414566 59304 414572 59316
rect 414624 59304 414630 59356
rect 59722 59236 59728 59288
rect 59780 59276 59786 59288
rect 94498 59276 94504 59288
rect 59780 59248 94504 59276
rect 59780 59236 59786 59248
rect 94498 59236 94504 59248
rect 94556 59236 94562 59288
rect 379606 59236 379612 59288
rect 379664 59276 379670 59288
rect 418154 59276 418160 59288
rect 379664 59248 418160 59276
rect 379664 59236 379670 59248
rect 418154 59236 418160 59248
rect 418212 59236 418218 59288
rect 57054 59168 57060 59220
rect 57112 59208 57118 59220
rect 95878 59208 95884 59220
rect 57112 59180 95884 59208
rect 57112 59168 57118 59180
rect 95878 59168 95884 59180
rect 95936 59168 95942 59220
rect 214650 59168 214656 59220
rect 214708 59208 214714 59220
rect 259454 59208 259460 59220
rect 214708 59180 259460 59208
rect 214708 59168 214714 59180
rect 259454 59168 259460 59180
rect 259512 59168 259518 59220
rect 371878 59168 371884 59220
rect 371936 59208 371942 59220
rect 410702 59208 410708 59220
rect 371936 59180 410708 59208
rect 371936 59168 371942 59180
rect 410702 59168 410708 59180
rect 410760 59168 410766 59220
rect 56502 59100 56508 59152
rect 56560 59140 56566 59152
rect 96982 59140 96988 59152
rect 56560 59112 96988 59140
rect 56560 59100 56566 59112
rect 96982 59100 96988 59112
rect 97040 59100 97046 59152
rect 214742 59100 214748 59152
rect 214800 59140 214806 59152
rect 261662 59140 261668 59152
rect 214800 59112 261668 59140
rect 214800 59100 214806 59112
rect 261662 59100 261668 59112
rect 261720 59100 261726 59152
rect 279234 59100 279240 59152
rect 279292 59140 279298 59152
rect 356606 59140 356612 59152
rect 279292 59112 356612 59140
rect 279292 59100 279298 59112
rect 356606 59100 356612 59112
rect 356664 59100 356670 59152
rect 376294 59100 376300 59152
rect 376352 59140 376358 59152
rect 419350 59140 419356 59152
rect 376352 59112 419356 59140
rect 376352 59100 376358 59112
rect 419350 59100 419356 59112
rect 419408 59100 419414 59152
rect 55030 59032 55036 59084
rect 55088 59072 55094 59084
rect 98086 59072 98092 59084
rect 55088 59044 98092 59072
rect 55088 59032 55094 59044
rect 98086 59032 98092 59044
rect 98144 59032 98150 59084
rect 205542 59032 205548 59084
rect 205600 59072 205606 59084
rect 290918 59072 290924 59084
rect 205600 59044 290924 59072
rect 205600 59032 205606 59044
rect 290918 59032 290924 59044
rect 290976 59032 290982 59084
rect 376478 59032 376484 59084
rect 376536 59072 376542 59084
rect 420638 59072 420644 59084
rect 376536 59044 420644 59072
rect 376536 59032 376542 59044
rect 420638 59032 420644 59044
rect 420696 59032 420702 59084
rect 56318 58964 56324 59016
rect 56376 59004 56382 59016
rect 102778 59004 102784 59016
rect 56376 58976 102784 59004
rect 56376 58964 56382 58976
rect 102778 58964 102784 58976
rect 102836 58964 102842 59016
rect 213822 58964 213828 59016
rect 213880 59004 213886 59016
rect 300854 59004 300860 59016
rect 213880 58976 300860 59004
rect 213880 58964 213886 58976
rect 300854 58964 300860 58976
rect 300912 58964 300918 59016
rect 376202 58964 376208 59016
rect 376260 59004 376266 59016
rect 421742 59004 421748 59016
rect 376260 58976 421748 59004
rect 376260 58964 376266 58976
rect 421742 58964 421748 58976
rect 421800 58964 421806 59016
rect 55858 58896 55864 58948
rect 55916 58936 55922 58948
rect 103882 58936 103888 58948
rect 55916 58908 103888 58936
rect 55916 58896 55922 58908
rect 103882 58896 103888 58908
rect 103940 58896 103946 58948
rect 212442 58896 212448 58948
rect 212500 58936 212506 58948
rect 315850 58936 315856 58948
rect 212500 58908 315856 58936
rect 212500 58896 212506 58908
rect 315850 58896 315856 58908
rect 315908 58896 315914 58948
rect 360838 58896 360844 58948
rect 360896 58936 360902 58948
rect 416038 58936 416044 58948
rect 360896 58908 416044 58936
rect 360896 58896 360902 58908
rect 416038 58896 416044 58908
rect 416096 58896 416102 58948
rect 59814 58828 59820 58880
rect 59872 58868 59878 58880
rect 108666 58868 108672 58880
rect 59872 58840 108672 58868
rect 59872 58828 59878 58840
rect 108666 58828 108672 58840
rect 108724 58828 108730 58880
rect 202782 58828 202788 58880
rect 202840 58868 202846 58880
rect 308490 58868 308496 58880
rect 202840 58840 308496 58868
rect 202840 58828 202846 58840
rect 308490 58828 308496 58840
rect 308548 58828 308554 58880
rect 358170 58828 358176 58880
rect 358228 58868 358234 58880
rect 423490 58868 423496 58880
rect 358228 58840 423496 58868
rect 358228 58828 358234 58840
rect 423490 58828 423496 58840
rect 423548 58828 423554 58880
rect 49602 58760 49608 58812
rect 49660 58800 49666 58812
rect 110966 58800 110972 58812
rect 49660 58772 110972 58800
rect 49660 58760 49666 58772
rect 110966 58760 110972 58772
rect 111024 58760 111030 58812
rect 209590 58760 209596 58812
rect 209648 58800 209654 58812
rect 320910 58800 320916 58812
rect 209648 58772 320916 58800
rect 209648 58760 209654 58772
rect 320910 58760 320916 58772
rect 320968 58760 320974 58812
rect 366450 58760 366456 58812
rect 366508 58800 366514 58812
rect 468478 58800 468484 58812
rect 366508 58772 468484 58800
rect 366508 58760 366514 58772
rect 468478 58760 468484 58772
rect 468536 58760 468542 58812
rect 50982 58692 50988 58744
rect 51040 58732 51046 58744
rect 148502 58732 148508 58744
rect 51040 58704 148508 58732
rect 51040 58692 51046 58704
rect 148502 58692 148508 58704
rect 148560 58692 148566 58744
rect 209498 58692 209504 58744
rect 209556 58732 209562 58744
rect 325878 58732 325884 58744
rect 209556 58704 325884 58732
rect 209556 58692 209562 58704
rect 325878 58692 325884 58704
rect 325936 58692 325942 58744
rect 363598 58692 363604 58744
rect 363656 58732 363662 58744
rect 475838 58732 475844 58744
rect 363656 58704 475844 58732
rect 363656 58692 363662 58704
rect 475838 58692 475844 58704
rect 475896 58692 475902 58744
rect 53006 58624 53012 58676
rect 53064 58664 53070 58676
rect 150894 58664 150900 58676
rect 53064 58636 150900 58664
rect 53064 58624 53070 58636
rect 150894 58624 150900 58636
rect 150952 58624 150958 58676
rect 219066 58624 219072 58676
rect 219124 58664 219130 58676
rect 428182 58664 428188 58676
rect 219124 58636 428188 58664
rect 219124 58624 219130 58636
rect 428182 58624 428188 58636
rect 428240 58624 428246 58676
rect 216398 58556 216404 58608
rect 216456 58596 216462 58608
rect 260650 58596 260656 58608
rect 216456 58568 260656 58596
rect 216456 58556 216462 58568
rect 260650 58556 260656 58568
rect 260708 58556 260714 58608
rect 375926 58556 375932 58608
rect 375984 58596 375990 58608
rect 404170 58596 404176 58608
rect 375984 58568 404176 58596
rect 375984 58556 375990 58568
rect 404170 58556 404176 58568
rect 404228 58556 404234 58608
rect 57882 57876 57888 57928
rect 57940 57916 57946 57928
rect 204898 57916 204904 57928
rect 57940 57888 204904 57916
rect 57940 57876 57946 57888
rect 204898 57876 204904 57888
rect 204956 57876 204962 57928
rect 211062 57876 211068 57928
rect 211120 57916 211126 57928
rect 323302 57916 323308 57928
rect 211120 57888 323308 57916
rect 211120 57876 211126 57888
rect 323302 57876 323308 57888
rect 323360 57876 323366 57928
rect 343174 57876 343180 57928
rect 343232 57916 343238 57928
rect 357526 57916 357532 57928
rect 343232 57888 357532 57916
rect 343232 57876 343238 57888
rect 357526 57876 357532 57888
rect 357584 57876 357590 57928
rect 376662 57876 376668 57928
rect 376720 57916 376726 57928
rect 485958 57916 485964 57928
rect 376720 57888 485964 57916
rect 376720 57876 376726 57888
rect 485958 57876 485964 57888
rect 486016 57876 486022 57928
rect 503254 57876 503260 57928
rect 503312 57916 503318 57928
rect 517606 57916 517612 57928
rect 503312 57888 517612 57916
rect 503312 57876 503318 57888
rect 517606 57876 517612 57888
rect 517664 57876 517670 57928
rect 51626 57808 51632 57860
rect 51684 57848 51690 57860
rect 145558 57848 145564 57860
rect 51684 57820 145564 57848
rect 51684 57808 51690 57820
rect 145558 57808 145564 57820
rect 145616 57808 145622 57860
rect 183278 57808 183284 57860
rect 183336 57848 183342 57860
rect 197446 57848 197452 57860
rect 183336 57820 197452 57848
rect 183336 57808 183342 57820
rect 197446 57808 197452 57820
rect 197504 57808 197510 57860
rect 206186 57808 206192 57860
rect 206244 57848 206250 57860
rect 313366 57848 313372 57860
rect 206244 57820 313372 57848
rect 206244 57808 206250 57820
rect 313366 57808 313372 57820
rect 313424 57808 313430 57860
rect 343450 57808 343456 57860
rect 343508 57848 343514 57860
rect 356698 57848 356704 57860
rect 343508 57820 356704 57848
rect 343508 57808 343514 57820
rect 356698 57808 356704 57820
rect 356756 57808 356762 57860
rect 365622 57808 365628 57860
rect 365680 57848 365686 57860
rect 470870 57848 470876 57860
rect 365680 57820 470876 57848
rect 365680 57808 365686 57820
rect 470870 57808 470876 57820
rect 470928 57808 470934 57860
rect 503530 57808 503536 57860
rect 503588 57848 503594 57860
rect 517882 57848 517888 57860
rect 503588 57820 517888 57848
rect 503588 57808 503594 57820
rect 517882 57808 517888 57820
rect 517940 57808 517946 57860
rect 43990 57740 43996 57792
rect 44048 57780 44054 57792
rect 123478 57780 123484 57792
rect 44048 57752 123484 57780
rect 44048 57740 44054 57752
rect 123478 57740 123484 57752
rect 123536 57740 123542 57792
rect 183462 57740 183468 57792
rect 183520 57780 183526 57792
rect 197354 57780 197360 57792
rect 183520 57752 197360 57780
rect 183520 57740 183526 57752
rect 197354 57740 197360 57752
rect 197412 57740 197418 57792
rect 218238 57740 218244 57792
rect 218296 57780 218302 57792
rect 318242 57780 318248 57792
rect 218296 57752 318248 57780
rect 218296 57740 218302 57752
rect 318242 57740 318248 57752
rect 318300 57740 318306 57792
rect 379422 57740 379428 57792
rect 379480 57780 379486 57792
rect 478414 57780 478420 57792
rect 379480 57752 478420 57780
rect 379480 57740 379486 57752
rect 478414 57740 478420 57752
rect 478472 57740 478478 57792
rect 53742 57672 53748 57724
rect 53800 57712 53806 57724
rect 133414 57712 133420 57724
rect 53800 57684 133420 57712
rect 53800 57672 53806 57684
rect 133414 57672 133420 57684
rect 133472 57672 133478 57724
rect 215110 57672 215116 57724
rect 215168 57712 215174 57724
rect 310974 57712 310980 57724
rect 215168 57684 310980 57712
rect 215168 57672 215174 57684
rect 310974 57672 310980 57684
rect 311032 57672 311038 57724
rect 367738 57672 367744 57724
rect 367796 57712 367802 57724
rect 465902 57712 465908 57724
rect 367796 57684 465908 57712
rect 367796 57672 367802 57684
rect 465902 57672 465908 57684
rect 465960 57672 465966 57724
rect 52362 57604 52368 57656
rect 52420 57644 52426 57656
rect 130838 57644 130844 57656
rect 52420 57616 130844 57644
rect 52420 57604 52426 57616
rect 130838 57604 130844 57616
rect 130896 57604 130902 57656
rect 208670 57604 208676 57656
rect 208728 57644 208734 57656
rect 303430 57644 303436 57656
rect 208728 57616 303436 57644
rect 208728 57604 208734 57616
rect 303430 57604 303436 57616
rect 303488 57604 303494 57656
rect 371142 57604 371148 57656
rect 371200 57644 371206 57656
rect 460934 57644 460940 57656
rect 371200 57616 460940 57644
rect 371200 57604 371206 57616
rect 460934 57604 460940 57616
rect 460992 57604 460998 57656
rect 54202 57536 54208 57588
rect 54260 57576 54266 57588
rect 128354 57576 128360 57588
rect 54260 57548 128360 57576
rect 54260 57536 54266 57548
rect 128354 57536 128360 57548
rect 128412 57536 128418 57588
rect 215662 57536 215668 57588
rect 215720 57576 215726 57588
rect 305822 57576 305828 57588
rect 215720 57548 305828 57576
rect 215720 57536 215726 57548
rect 305822 57536 305828 57548
rect 305880 57536 305886 57588
rect 369118 57536 369124 57588
rect 369176 57576 369182 57588
rect 445846 57576 445852 57588
rect 369176 57548 445852 57576
rect 369176 57536 369182 57548
rect 445846 57536 445852 57548
rect 445904 57536 445910 57588
rect 44082 57468 44088 57520
rect 44140 57508 44146 57520
rect 44140 57480 45554 57508
rect 44140 57468 44146 57480
rect 45526 57440 45554 57480
rect 57238 57468 57244 57520
rect 57296 57508 57302 57520
rect 57882 57508 57888 57520
rect 57296 57480 57888 57508
rect 57296 57468 57302 57480
rect 57882 57468 57888 57480
rect 57940 57468 57946 57520
rect 115934 57508 115940 57520
rect 58820 57480 115940 57508
rect 58820 57440 58848 57480
rect 115934 57468 115940 57480
rect 115992 57468 115998 57520
rect 210970 57468 210976 57520
rect 211028 57508 211034 57520
rect 295886 57508 295892 57520
rect 211028 57480 295892 57508
rect 211028 57468 211034 57480
rect 295886 57468 295892 57480
rect 295944 57468 295950 57520
rect 362218 57468 362224 57520
rect 362276 57508 362282 57520
rect 438486 57508 438492 57520
rect 362276 57480 438492 57508
rect 362276 57468 362282 57480
rect 438486 57468 438492 57480
rect 438544 57468 438550 57520
rect 45526 57412 58848 57440
rect 59998 57400 60004 57452
rect 60056 57440 60062 57452
rect 125870 57440 125876 57452
rect 60056 57412 125876 57440
rect 60056 57400 60062 57412
rect 125870 57400 125876 57412
rect 125928 57400 125934 57452
rect 210418 57400 210424 57452
rect 210476 57440 210482 57452
rect 293310 57440 293316 57452
rect 210476 57412 293316 57440
rect 210476 57400 210482 57412
rect 293310 57400 293316 57412
rect 293368 57400 293374 57452
rect 364978 57400 364984 57452
rect 365036 57440 365042 57452
rect 433518 57440 433524 57452
rect 365036 57412 433524 57440
rect 365036 57400 365042 57412
rect 433518 57400 433524 57412
rect 433576 57400 433582 57452
rect 55950 57332 55956 57384
rect 56008 57372 56014 57384
rect 99374 57372 99380 57384
rect 56008 57344 99380 57372
rect 56008 57332 56014 57344
rect 99374 57332 99380 57344
rect 99432 57332 99438 57384
rect 218790 57332 218796 57384
rect 218848 57372 218854 57384
rect 298094 57372 298100 57384
rect 218848 57344 298100 57372
rect 218848 57332 218854 57344
rect 298094 57332 298100 57344
rect 298152 57332 298158 57384
rect 371970 57332 371976 57384
rect 372028 57372 372034 57384
rect 435910 57372 435916 57384
rect 372028 57344 435916 57372
rect 372028 57332 372034 57344
rect 435910 57332 435916 57344
rect 435968 57332 435974 57384
rect 59262 57264 59268 57316
rect 59320 57304 59326 57316
rect 93578 57304 93584 57316
rect 59320 57276 93584 57304
rect 59320 57264 59326 57276
rect 93578 57264 93584 57276
rect 93636 57264 93642 57316
rect 215202 57264 215208 57316
rect 215260 57304 215266 57316
rect 287606 57304 287612 57316
rect 215260 57276 287612 57304
rect 215260 57264 215266 57276
rect 287606 57264 287612 57276
rect 287664 57264 287670 57316
rect 370498 57264 370504 57316
rect 370556 57304 370562 57316
rect 430942 57304 430948 57316
rect 370556 57276 430948 57304
rect 370556 57264 370562 57276
rect 430942 57264 430948 57276
rect 431000 57264 431006 57316
rect 51718 57196 51724 57248
rect 51776 57236 51782 57248
rect 78214 57236 78220 57248
rect 51776 57208 78220 57236
rect 51776 57196 51782 57208
rect 78214 57196 78220 57208
rect 78272 57196 78278 57248
rect 218698 57196 218704 57248
rect 218756 57236 218762 57248
rect 258350 57236 258356 57248
rect 218756 57208 258356 57236
rect 218756 57196 218762 57208
rect 258350 57196 258356 57208
rect 258408 57196 258414 57248
rect 378410 57196 378416 57248
rect 378468 57236 378474 57248
rect 415486 57236 415492 57248
rect 378468 57208 415492 57236
rect 378468 57196 378474 57208
rect 415486 57196 415492 57208
rect 415544 57196 415550 57248
rect 54754 57128 54760 57180
rect 54812 57168 54818 57180
rect 76006 57168 76012 57180
rect 54812 57140 76012 57168
rect 54812 57128 54818 57140
rect 76006 57128 76012 57140
rect 76064 57128 76070 57180
rect 54294 56516 54300 56568
rect 54352 56556 54358 56568
rect 116670 56556 116676 56568
rect 54352 56528 116676 56556
rect 54352 56516 54358 56528
rect 116670 56516 116676 56528
rect 116728 56516 116734 56568
rect 219986 56516 219992 56568
rect 220044 56556 220050 56568
rect 408310 56556 408316 56568
rect 220044 56528 408316 56556
rect 220044 56516 220050 56528
rect 408310 56516 408316 56528
rect 408368 56516 408374 56568
rect 53098 56448 53104 56500
rect 53156 56488 53162 56500
rect 113818 56488 113824 56500
rect 53156 56460 113824 56488
rect 53156 56448 53162 56460
rect 113818 56448 113824 56460
rect 113876 56448 113882 56500
rect 213546 56448 213552 56500
rect 213604 56488 213610 56500
rect 273254 56488 273260 56500
rect 213604 56460 273260 56488
rect 213604 56448 213610 56460
rect 273254 56448 273260 56460
rect 273312 56448 273318 56500
rect 376570 56448 376576 56500
rect 376628 56488 376634 56500
rect 436370 56488 436376 56500
rect 376628 56460 436376 56488
rect 376628 56448 376634 56460
rect 436370 56448 436376 56460
rect 436428 56448 436434 56500
rect 52086 56380 52092 56432
rect 52144 56420 52150 56432
rect 112070 56420 112076 56432
rect 52144 56392 112076 56420
rect 52144 56380 52150 56392
rect 112070 56380 112076 56392
rect 112128 56380 112134 56432
rect 216306 56380 216312 56432
rect 216364 56420 216370 56432
rect 276934 56420 276940 56432
rect 216364 56392 276940 56420
rect 216364 56380 216370 56392
rect 276934 56380 276940 56392
rect 276992 56380 276998 56432
rect 375282 56380 375288 56432
rect 375340 56420 375346 56432
rect 434622 56420 434628 56432
rect 375340 56392 434628 56420
rect 375340 56380 375346 56392
rect 434622 56380 434628 56392
rect 434680 56380 434686 56432
rect 53650 56312 53656 56364
rect 53708 56352 53714 56364
rect 109494 56352 109500 56364
rect 53708 56324 109500 56352
rect 53708 56312 53714 56324
rect 109494 56312 109500 56324
rect 109552 56312 109558 56364
rect 215018 56312 215024 56364
rect 215076 56352 215082 56364
rect 271046 56352 271052 56364
rect 215076 56324 271052 56352
rect 215076 56312 215082 56324
rect 271046 56312 271052 56324
rect 271104 56312 271110 56364
rect 374914 56312 374920 56364
rect 374972 56352 374978 56364
rect 432230 56352 432236 56364
rect 374972 56324 432236 56352
rect 374972 56312 374978 56324
rect 432230 56312 432236 56324
rect 432288 56312 432294 56364
rect 42702 56244 42708 56296
rect 42760 56284 42766 56296
rect 90726 56284 90732 56296
rect 42760 56256 90732 56284
rect 42760 56244 42766 56256
rect 90726 56244 90732 56256
rect 90784 56244 90790 56296
rect 219894 56244 219900 56296
rect 219952 56284 219958 56296
rect 268470 56284 268476 56296
rect 219952 56256 268476 56284
rect 219952 56244 219958 56256
rect 268470 56244 268476 56256
rect 268528 56244 268534 56296
rect 379238 56244 379244 56296
rect 379296 56284 379302 56296
rect 412634 56284 412640 56296
rect 379296 56256 412640 56284
rect 379296 56244 379302 56256
rect 412634 56244 412640 56256
rect 412692 56244 412698 56296
rect 58618 56176 58624 56228
rect 58676 56216 58682 56228
rect 92198 56216 92204 56228
rect 58676 56188 92204 56216
rect 58676 56176 58682 56188
rect 92198 56176 92204 56188
rect 92256 56176 92262 56228
rect 218606 56176 218612 56228
rect 218664 56216 218670 56228
rect 266354 56216 266360 56228
rect 218664 56188 266360 56216
rect 218664 56176 218670 56188
rect 266354 56176 266360 56188
rect 266412 56176 266418 56228
rect 376386 56176 376392 56228
rect 376444 56216 376450 56228
rect 408678 56216 408684 56228
rect 376444 56188 408684 56216
rect 376444 56176 376450 56188
rect 408678 56176 408684 56188
rect 408736 56176 408742 56228
rect 56410 56108 56416 56160
rect 56468 56148 56474 56160
rect 88702 56148 88708 56160
rect 56468 56120 88708 56148
rect 56468 56108 56474 56120
rect 88702 56108 88708 56120
rect 88760 56108 88766 56160
rect 215754 56108 215760 56160
rect 215812 56148 215818 56160
rect 250070 56148 250076 56160
rect 215812 56120 250076 56148
rect 215812 56108 215818 56120
rect 250070 56108 250076 56120
rect 250128 56108 250134 56160
rect 379330 56108 379336 56160
rect 379388 56148 379394 56160
rect 411254 56148 411260 56160
rect 379388 56120 411260 56148
rect 379388 56108 379394 56120
rect 411254 56108 411260 56120
rect 411312 56108 411318 56160
rect 54846 56040 54852 56092
rect 54904 56080 54910 56092
rect 86494 56080 86500 56092
rect 54904 56052 86500 56080
rect 54904 56040 54910 56052
rect 86494 56040 86500 56052
rect 86552 56040 86558 56092
rect 217042 56040 217048 56092
rect 217100 56080 217106 56092
rect 251910 56080 251916 56092
rect 217100 56052 251916 56080
rect 217100 56040 217106 56052
rect 251910 56040 251916 56052
rect 251968 56040 251974 56092
rect 373810 56040 373816 56092
rect 373868 56080 373874 56092
rect 401686 56080 401692 56092
rect 373868 56052 401692 56080
rect 373868 56040 373874 56052
rect 401686 56040 401692 56052
rect 401744 56040 401750 56092
rect 51994 55972 52000 56024
rect 52052 56012 52058 56024
rect 81894 56012 81900 56024
rect 52052 55984 81900 56012
rect 52052 55972 52058 55984
rect 81894 55972 81900 55984
rect 81952 55972 81958 56024
rect 216122 55972 216128 56024
rect 216180 56012 216186 56024
rect 247678 56012 247684 56024
rect 216180 55984 247684 56012
rect 216180 55972 216186 55984
rect 247678 55972 247684 55984
rect 247736 55972 247742 56024
rect 374730 55972 374736 56024
rect 374788 56012 374794 56024
rect 399478 56012 399484 56024
rect 374788 55984 399484 56012
rect 374788 55972 374794 55984
rect 399478 55972 399484 55984
rect 399536 55972 399542 56024
rect 58710 55904 58716 55956
rect 58768 55944 58774 55956
rect 85390 55944 85396 55956
rect 58768 55916 85396 55944
rect 58768 55904 58774 55916
rect 85390 55904 85396 55916
rect 85448 55904 85454 55956
rect 216030 55904 216036 55956
rect 216088 55944 216094 55956
rect 245286 55944 245292 55956
rect 216088 55916 245292 55944
rect 216088 55904 216094 55916
rect 245286 55904 245292 55916
rect 245344 55904 245350 55956
rect 53466 55836 53472 55888
rect 53524 55876 53530 55888
rect 79502 55876 79508 55888
rect 53524 55848 79508 55876
rect 53524 55836 53530 55848
rect 79502 55836 79508 55848
rect 79560 55836 79566 55888
rect 213270 55836 213276 55888
rect 213328 55876 213334 55888
rect 239214 55876 239220 55888
rect 213328 55848 239220 55876
rect 213328 55836 213334 55848
rect 239214 55836 239220 55848
rect 239272 55836 239278 55888
rect 213178 55768 213184 55820
rect 213236 55808 213242 55820
rect 241606 55808 241612 55820
rect 213236 55780 241612 55808
rect 213236 55768 213242 55780
rect 241606 55768 241612 55780
rect 241664 55768 241670 55820
rect 50890 55156 50896 55208
rect 50948 55196 50954 55208
rect 114554 55196 114560 55208
rect 50948 55168 114560 55196
rect 50948 55156 50954 55168
rect 114554 55156 114560 55168
rect 114612 55156 114618 55208
rect 218882 55156 218888 55208
rect 218940 55196 218946 55208
rect 245654 55196 245660 55208
rect 218940 55168 245660 55196
rect 218940 55156 218946 55168
rect 245654 55156 245660 55168
rect 245712 55156 245718 55208
rect 378778 55156 378784 55208
rect 378836 55196 378842 55208
rect 407206 55196 407212 55208
rect 378836 55168 407212 55196
rect 378836 55156 378842 55168
rect 407206 55156 407212 55168
rect 407264 55156 407270 55208
rect 53558 55088 53564 55140
rect 53616 55128 53622 55140
rect 113266 55128 113272 55140
rect 53616 55100 113272 55128
rect 53616 55088 53622 55100
rect 113266 55088 113272 55100
rect 113324 55088 113330 55140
rect 215938 55088 215944 55140
rect 215996 55128 216002 55140
rect 271874 55128 271880 55140
rect 215996 55100 271880 55128
rect 215996 55088 216002 55100
rect 271874 55088 271880 55100
rect 271932 55088 271938 55140
rect 379054 55088 379060 55140
rect 379112 55128 379118 55140
rect 437474 55128 437480 55140
rect 379112 55100 437480 55128
rect 379112 55088 379118 55100
rect 437474 55088 437480 55100
rect 437532 55088 437538 55140
rect 52178 55020 52184 55072
rect 52236 55060 52242 55072
rect 110414 55060 110420 55072
rect 52236 55032 110420 55060
rect 52236 55020 52242 55032
rect 110414 55020 110420 55032
rect 110472 55020 110478 55072
rect 219526 55020 219532 55072
rect 219584 55060 219590 55072
rect 266446 55060 266452 55072
rect 219584 55032 266452 55060
rect 219584 55020 219590 55032
rect 266446 55020 266452 55032
rect 266504 55020 266510 55072
rect 375190 55020 375196 55072
rect 375248 55060 375254 55072
rect 433426 55060 433432 55072
rect 375248 55032 433432 55060
rect 375248 55020 375254 55032
rect 433426 55020 433432 55032
rect 433484 55020 433490 55072
rect 59906 54952 59912 55004
rect 59964 54992 59970 55004
rect 106274 54992 106280 55004
rect 59964 54964 106280 54992
rect 59964 54952 59970 54964
rect 106274 54952 106280 54964
rect 106332 54952 106338 55004
rect 219618 54952 219624 55004
rect 219676 54992 219682 55004
rect 264974 54992 264980 55004
rect 219676 54964 264980 54992
rect 219676 54952 219682 54964
rect 264974 54952 264980 54964
rect 265032 54952 265038 55004
rect 375006 54952 375012 55004
rect 375064 54992 375070 55004
rect 430574 54992 430580 55004
rect 375064 54964 430580 54992
rect 375064 54952 375070 54964
rect 430574 54952 430580 54964
rect 430632 54952 430638 55004
rect 56962 54884 56968 54936
rect 57020 54924 57026 54936
rect 91186 54924 91192 54936
rect 57020 54896 91192 54924
rect 57020 54884 57026 54896
rect 91186 54884 91192 54896
rect 91244 54884 91250 54936
rect 218330 54884 218336 54936
rect 218388 54924 218394 54936
rect 263594 54924 263600 54936
rect 218388 54896 263600 54924
rect 218388 54884 218394 54896
rect 263594 54884 263600 54896
rect 263652 54884 263658 54936
rect 375098 54884 375104 54936
rect 375156 54924 375162 54936
rect 429194 54924 429200 54936
rect 375156 54896 429200 54924
rect 375156 54884 375162 54896
rect 429194 54884 429200 54896
rect 429252 54884 429258 54936
rect 53190 54816 53196 54868
rect 53248 54856 53254 54868
rect 86954 54856 86960 54868
rect 53248 54828 86960 54856
rect 53248 54816 53254 54828
rect 86954 54816 86960 54828
rect 87012 54816 87018 54868
rect 219710 54816 219716 54868
rect 219768 54856 219774 54868
rect 253934 54856 253940 54868
rect 219768 54828 253940 54856
rect 219768 54816 219774 54828
rect 253934 54816 253940 54828
rect 253992 54816 253998 54868
rect 379790 54816 379796 54868
rect 379848 54856 379854 54868
rect 426434 54856 426440 54868
rect 379848 54828 426440 54856
rect 379848 54816 379854 54828
rect 426434 54816 426440 54828
rect 426492 54816 426498 54868
rect 59078 54748 59084 54800
rect 59136 54788 59142 54800
rect 92474 54788 92480 54800
rect 59136 54760 92480 54788
rect 59136 54748 59142 54760
rect 92474 54748 92480 54760
rect 92532 54748 92538 54800
rect 218422 54748 218428 54800
rect 218480 54788 218486 54800
rect 252554 54788 252560 54800
rect 218480 54760 252560 54788
rect 218480 54748 218486 54760
rect 252554 54748 252560 54760
rect 252612 54748 252618 54800
rect 379514 54748 379520 54800
rect 379572 54788 379578 54800
rect 426526 54788 426532 54800
rect 379572 54760 426532 54788
rect 379572 54748 379578 54760
rect 426526 54748 426532 54760
rect 426584 54748 426590 54800
rect 59170 54680 59176 54732
rect 59228 54720 59234 54732
rect 89806 54720 89812 54732
rect 59228 54692 89812 54720
rect 59228 54680 59234 54692
rect 89806 54680 89812 54692
rect 89864 54680 89870 54732
rect 219250 54680 219256 54732
rect 219308 54720 219314 54732
rect 251174 54720 251180 54732
rect 219308 54692 251180 54720
rect 219308 54680 219314 54692
rect 251174 54680 251180 54692
rect 251232 54680 251238 54732
rect 377582 54680 377588 54732
rect 377640 54720 377646 54732
rect 411346 54720 411352 54732
rect 377640 54692 411352 54720
rect 377640 54680 377646 54692
rect 411346 54680 411352 54692
rect 411404 54680 411410 54732
rect 54938 54612 54944 54664
rect 54996 54652 55002 54664
rect 80054 54652 80060 54664
rect 54996 54624 80060 54652
rect 54996 54612 55002 54624
rect 80054 54612 80060 54624
rect 80112 54612 80118 54664
rect 217134 54612 217140 54664
rect 217192 54652 217198 54664
rect 248414 54652 248420 54664
rect 217192 54624 248420 54652
rect 217192 54612 217198 54624
rect 248414 54612 248420 54624
rect 248472 54612 248478 54664
rect 378042 54612 378048 54664
rect 378100 54652 378106 54664
rect 409874 54652 409880 54664
rect 378100 54624 409880 54652
rect 378100 54612 378106 54624
rect 409874 54612 409880 54624
rect 409932 54612 409938 54664
rect 214834 54544 214840 54596
rect 214892 54584 214898 54596
rect 244366 54584 244372 54596
rect 214892 54556 244372 54584
rect 214892 54544 214898 54556
rect 244366 54544 244372 54556
rect 244424 54544 244430 54596
rect 376018 54544 376024 54596
rect 376076 54584 376082 54596
rect 405826 54584 405832 54596
rect 376076 54556 405832 54584
rect 376076 54544 376082 54556
rect 405826 54544 405832 54556
rect 405884 54544 405890 54596
rect 216490 54476 216496 54528
rect 216548 54516 216554 54528
rect 242894 54516 242900 54528
rect 216548 54488 242900 54516
rect 216548 54476 216554 54488
rect 242894 54476 242900 54488
rect 242952 54476 242958 54528
rect 374822 54476 374828 54528
rect 374880 54516 374886 54528
rect 404354 54516 404360 54528
rect 374880 54488 404360 54516
rect 374880 54476 374886 54488
rect 404354 54476 404360 54488
rect 404412 54476 404418 54528
rect 213362 54408 213368 54460
rect 213420 54448 213426 54460
rect 273346 54448 273352 54460
rect 213420 54420 273352 54448
rect 213420 54408 213426 54420
rect 273346 54408 273352 54420
rect 273404 54408 273410 54460
rect 372522 54408 372528 54460
rect 372580 54448 372586 54460
rect 434714 54448 434720 54460
rect 372580 54420 434720 54448
rect 372580 54408 372586 54420
rect 434714 54408 434720 54420
rect 434772 54408 434778 54460
rect 213454 54340 213460 54392
rect 213512 54380 213518 54392
rect 237374 54380 237380 54392
rect 213512 54352 237380 54380
rect 213512 54340 213518 54352
rect 237374 54340 237380 54352
rect 237432 54340 237438 54392
rect 374638 54340 374644 54392
rect 374696 54380 374702 54392
rect 397454 54380 397460 54392
rect 374696 54352 397460 54380
rect 374696 54340 374702 54352
rect 397454 54340 397460 54352
rect 397512 54340 397518 54392
rect 214558 54272 214564 54324
rect 214616 54312 214622 54324
rect 240134 54312 240140 54324
rect 214616 54284 240140 54312
rect 214616 54272 214622 54284
rect 240134 54272 240140 54284
rect 240192 54272 240198 54324
rect 372430 54272 372436 54324
rect 372488 54312 372494 54324
rect 400214 54312 400220 54324
rect 372488 54284 400220 54312
rect 372488 54272 372494 54284
rect 400214 54272 400220 54284
rect 400272 54272 400278 54324
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 10318 20652 10324 20664
rect 3476 20624 10324 20652
rect 3476 20612 3482 20624
rect 10318 20612 10324 20624
rect 10376 20612 10382 20664
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 57238 3448 57244 3460
rect 624 3420 57244 3448
rect 624 3408 630 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 125870 3408 125876 3460
rect 125928 3448 125934 3460
rect 366358 3448 366364 3460
rect 125928 3420 366364 3448
rect 125928 3408 125934 3420
rect 366358 3408 366364 3420
rect 366416 3408 366422 3460
<< via1 >>
rect 235172 700408 235224 700460
rect 305644 700408 305696 700460
rect 429844 700408 429896 700460
rect 434720 700408 434772 700460
rect 170312 700340 170364 700392
rect 434904 700340 434956 700392
rect 57796 700272 57848 700324
rect 543464 700272 543516 700324
rect 147588 683136 147640 683188
rect 580172 683136 580224 683188
rect 299480 640976 299532 641028
rect 405740 640976 405792 641028
rect 104900 639548 104952 639600
rect 434812 639548 434864 639600
rect 3424 638188 3476 638240
rect 318156 638188 318208 638240
rect 364340 638188 364392 638240
rect 428280 638188 428332 638240
rect 40040 636828 40092 636880
rect 320824 636828 320876 636880
rect 307024 635740 307076 635792
rect 355600 635740 355652 635792
rect 322480 635672 322532 635724
rect 346584 635672 346636 635724
rect 322296 635604 322348 635656
rect 432880 635604 432932 635656
rect 318064 635536 318116 635588
rect 392308 635536 392360 635588
rect 323952 635468 324004 635520
rect 369124 635468 369176 635520
rect 319444 635400 319496 635452
rect 364616 635400 364668 635452
rect 316776 635332 316828 635384
rect 342260 635332 342312 635384
rect 361396 635332 361448 635384
rect 414848 635332 414900 635384
rect 324872 635264 324924 635316
rect 378140 635264 378192 635316
rect 353300 635196 353352 635248
rect 410340 635196 410392 635248
rect 313924 635128 313976 635180
rect 374000 635128 374052 635180
rect 321008 635060 321060 635112
rect 387800 635060 387852 635112
rect 314016 634992 314068 635044
rect 383660 634992 383712 635044
rect 323860 634924 323912 634976
rect 401600 634924 401652 634976
rect 322388 634856 322440 634908
rect 337568 634856 337620 634908
rect 323768 634788 323820 634840
rect 328644 634788 328696 634840
rect 391940 634788 391992 634840
rect 420000 634788 420052 634840
rect 457444 634788 457496 634840
rect 323676 634312 323728 634364
rect 436192 634312 436244 634364
rect 322572 634244 322624 634296
rect 436100 634244 436152 634296
rect 236644 634176 236696 634228
rect 360200 634176 360252 634228
rect 144920 634108 144972 634160
rect 145012 634040 145064 634092
rect 156604 634040 156656 634092
rect 239404 634108 239456 634160
rect 257068 634108 257120 634160
rect 322664 634108 322716 634160
rect 457720 634108 457772 634160
rect 207664 634040 207716 634092
rect 238208 634040 238260 634092
rect 251364 634040 251416 634092
rect 324228 634040 324280 634092
rect 494060 634040 494112 634092
rect 109960 633972 110012 634024
rect 120908 633972 120960 634024
rect 148876 633972 148928 634024
rect 172888 633972 172940 634024
rect 226340 633972 226392 634024
rect 300308 633972 300360 634024
rect 316960 633972 317012 634024
rect 457536 633972 457588 634024
rect 112536 633904 112588 633956
rect 122932 633904 122984 633956
rect 140780 633904 140832 633956
rect 167092 633904 167144 633956
rect 214012 633904 214064 633956
rect 289268 633904 289320 633956
rect 314200 633904 314252 633956
rect 456800 633904 456852 633956
rect 86776 633836 86828 633888
rect 124312 633836 124364 633888
rect 148784 633836 148836 633888
rect 176108 633836 176160 633888
rect 231124 633836 231176 633888
rect 248788 633836 248840 633888
rect 304264 633836 304316 633888
rect 457628 633836 457680 633888
rect 115664 633768 115716 633820
rect 124588 633768 124640 633820
rect 149796 633768 149848 633820
rect 190552 633768 190604 633820
rect 234620 633768 234672 633820
rect 396816 633768 396868 633820
rect 106648 633700 106700 633752
rect 121000 633700 121052 633752
rect 142160 633700 142212 633752
rect 184480 633700 184532 633752
rect 239588 633700 239640 633752
rect 274640 633700 274692 633752
rect 304356 633700 304408 633752
rect 471612 633700 471664 633752
rect 56508 633632 56560 633684
rect 77300 633632 77352 633684
rect 104072 633632 104124 633684
rect 122196 633632 122248 633684
rect 156604 633632 156656 633684
rect 196072 633632 196124 633684
rect 213920 633632 213972 633684
rect 245660 633632 245712 633684
rect 249340 633632 249392 633684
rect 295524 633632 295576 633684
rect 314108 633632 314160 633684
rect 483204 633632 483256 633684
rect 55036 633564 55088 633616
rect 80244 633564 80296 633616
rect 100668 633564 100720 633616
rect 124496 633564 124548 633616
rect 147496 633564 147548 633616
rect 199292 633564 199344 633616
rect 235264 633564 235316 633616
rect 291844 633564 291896 633616
rect 322204 633564 322256 633616
rect 494796 633564 494848 633616
rect 55128 633496 55180 633548
rect 91836 633496 91888 633548
rect 95056 633496 95108 633548
rect 121644 633496 121696 633548
rect 133880 633496 133932 633548
rect 149980 633496 150032 633548
rect 54852 633428 54904 633480
rect 88708 633428 88760 633480
rect 147404 633428 147456 633480
rect 149704 633428 149756 633480
rect 201868 633496 201920 633548
rect 205548 633496 205600 633548
rect 212632 633496 212684 633548
rect 237380 633496 237432 633548
rect 254492 633496 254544 633548
rect 320916 633496 320968 633548
rect 501236 633496 501288 633548
rect 164516 633428 164568 633480
rect 255320 633428 255372 633480
rect 262956 633428 263008 633480
rect 316868 633428 316920 633480
rect 512184 633428 512236 633480
rect 223580 632952 223632 633004
rect 249340 632952 249392 633004
rect 222200 632884 222252 632936
rect 255320 632884 255372 632936
rect 3516 632816 3568 632868
rect 353300 632816 353352 632868
rect 3608 632748 3660 632800
rect 361396 632748 361448 632800
rect 237840 632680 237892 632732
rect 391940 632680 391992 632732
rect 238944 632476 238996 632528
rect 580172 632476 580224 632528
rect 3424 632408 3476 632460
rect 323584 632408 323636 632460
rect 319628 632340 319680 632392
rect 436284 632340 436336 632392
rect 239036 632272 239088 632324
rect 433340 632272 433392 632324
rect 317052 632204 317104 632256
rect 512092 632204 512144 632256
rect 319536 632136 319588 632188
rect 512000 632136 512052 632188
rect 146116 631252 146168 631304
rect 155500 631252 155552 631304
rect 228364 631252 228416 631304
rect 280252 631252 280304 631304
rect 124864 631184 124916 631236
rect 187700 631184 187752 631236
rect 233884 631184 233936 631236
rect 266544 631184 266596 631236
rect 148968 631116 149020 631168
rect 158720 631116 158772 631168
rect 238116 631116 238168 631168
rect 277676 631116 277728 631168
rect 144184 631048 144236 631100
rect 161480 631048 161532 631100
rect 231216 631048 231268 631100
rect 271972 631048 272024 631100
rect 56416 630980 56468 631032
rect 65524 630980 65576 631032
rect 149888 630980 149940 631032
rect 170312 630980 170364 631032
rect 217324 630980 217376 631032
rect 260380 630980 260432 631032
rect 56324 630912 56376 630964
rect 71228 630912 71280 630964
rect 83464 630912 83516 630964
rect 124404 630912 124456 630964
rect 136640 630912 136692 630964
rect 178684 630912 178736 630964
rect 214564 630912 214616 630964
rect 268660 630912 268712 630964
rect 59360 630844 59412 630896
rect 97908 630844 97960 630896
rect 140044 630844 140096 630896
rect 193496 630844 193548 630896
rect 220176 630844 220228 630896
rect 283564 630844 283616 630896
rect 57704 630776 57756 630828
rect 74632 630776 74684 630828
rect 124220 630776 124272 630828
rect 182088 630776 182140 630828
rect 220084 630776 220136 630828
rect 286140 630776 286192 630828
rect 54944 630708 54996 630760
rect 62948 630708 63000 630760
rect 69296 630708 69348 630760
rect 125784 630708 125836 630760
rect 148324 630708 148376 630760
rect 153108 630708 153160 630760
rect 215944 630708 215996 630760
rect 297732 630708 297784 630760
rect 57888 630640 57940 630692
rect 146208 630640 146260 630692
rect 237840 630640 237892 630692
rect 239496 630640 239548 630692
rect 242900 630640 242952 630692
rect 118148 630368 118200 630420
rect 121460 630368 121512 630420
rect 215300 629892 215352 629944
rect 237380 629892 237432 629944
rect 144276 627920 144328 627972
rect 146300 627920 146352 627972
rect 217416 627920 217468 627972
rect 237380 627920 237432 627972
rect 465448 627920 465500 627972
rect 580264 627920 580316 627972
rect 238852 627784 238904 627836
rect 239772 627784 239824 627836
rect 309784 626560 309836 626612
rect 321560 626560 321612 626612
rect 233240 622412 233292 622464
rect 237380 622412 237432 622464
rect 311164 622412 311216 622464
rect 321560 622412 321612 622464
rect 140872 619624 140924 619676
rect 146300 619624 146352 619676
rect 232504 619624 232556 619676
rect 237380 619624 237432 619676
rect 316684 616836 316736 616888
rect 321560 616836 321612 616888
rect 132500 615476 132552 615528
rect 146300 615476 146352 615528
rect 222844 615476 222896 615528
rect 237380 615476 237432 615528
rect 223672 612756 223724 612808
rect 237380 612756 237432 612808
rect 312544 612756 312596 612808
rect 321560 612756 321612 612808
rect 218060 609968 218112 610020
rect 237380 609968 237432 610020
rect 312636 607180 312688 607232
rect 321560 607180 321612 607232
rect 307116 603100 307168 603152
rect 321560 603100 321612 603152
rect 229744 600312 229796 600364
rect 237380 600312 237432 600364
rect 129004 597524 129056 597576
rect 146300 597524 146352 597576
rect 217508 597524 217560 597576
rect 237380 597524 237432 597576
rect 307208 597524 307260 597576
rect 321560 597524 321612 597576
rect 302700 596776 302752 596828
rect 322664 596776 322716 596828
rect 124128 596164 124180 596216
rect 145564 596164 145616 596216
rect 214656 594804 214708 594856
rect 237380 594804 237432 594856
rect 57428 591336 57480 591388
rect 58624 591336 58676 591388
rect 220268 590656 220320 590708
rect 237380 590656 237432 590708
rect 305736 589296 305788 589348
rect 321560 589296 321612 589348
rect 231860 587868 231912 587920
rect 237380 587868 237432 587920
rect 125600 585148 125652 585200
rect 146300 585148 146352 585200
rect 235356 585148 235408 585200
rect 237380 585148 237432 585200
rect 307300 583720 307352 583772
rect 321560 583720 321612 583772
rect 130384 582360 130436 582412
rect 146300 582360 146352 582412
rect 57796 581612 57848 581664
rect 58716 581612 58768 581664
rect 139400 579640 139452 579692
rect 146300 579640 146352 579692
rect 216036 579640 216088 579692
rect 237380 579640 237432 579692
rect 317144 579640 317196 579692
rect 321560 579640 321612 579692
rect 513012 579640 513064 579692
rect 560944 579640 560996 579692
rect 226432 576852 226484 576904
rect 237380 576852 237432 576904
rect 311256 574064 311308 574116
rect 321560 574064 321612 574116
rect 218152 572704 218204 572756
rect 237380 572704 237432 572756
rect 220360 569916 220412 569968
rect 237380 569916 237432 569968
rect 318156 569848 318208 569900
rect 321560 569848 321612 569900
rect 57152 569168 57204 569220
rect 59912 569168 59964 569220
rect 3424 568488 3476 568540
rect 307300 568488 307352 568540
rect 57336 568420 57388 568472
rect 60740 568420 60792 568472
rect 113180 568420 113232 568472
rect 122288 568420 122340 568472
rect 145564 568420 145616 568472
rect 214104 568420 214156 568472
rect 302700 568420 302752 568472
rect 106280 568352 106332 568404
rect 124588 568352 124640 568404
rect 147128 568352 147180 568404
rect 151084 568352 151136 568404
rect 288532 568352 288584 568404
rect 316868 568352 316920 568404
rect 99564 568284 99616 568336
rect 123576 568284 123628 568336
rect 288624 568284 288676 568336
rect 316960 568284 317012 568336
rect 96712 568216 96764 568268
rect 122932 568216 122984 568268
rect 287060 568216 287112 568268
rect 317052 568216 317104 568268
rect 87052 568148 87104 568200
rect 121368 568148 121420 568200
rect 149704 568148 149756 568200
rect 154764 568148 154816 568200
rect 204904 568148 204956 568200
rect 212908 568148 212960 568200
rect 266360 568148 266412 568200
rect 314016 568148 314068 568200
rect 58808 568080 58860 568132
rect 67640 568080 67692 568132
rect 93860 568080 93912 568132
rect 124496 568080 124548 568132
rect 147496 568080 147548 568132
rect 156052 568080 156104 568132
rect 164424 568080 164476 568132
rect 212632 568080 212684 568132
rect 260840 568080 260892 568132
rect 319628 568080 319680 568132
rect 58992 568012 59044 568064
rect 74540 568012 74592 568064
rect 98092 568012 98144 568064
rect 120908 568012 120960 568064
rect 121460 568012 121512 568064
rect 211252 568012 211304 568064
rect 258080 568012 258132 568064
rect 322572 568012 322624 568064
rect 54852 567944 54904 567996
rect 78680 567944 78732 567996
rect 86960 567944 87012 567996
rect 121000 567944 121052 567996
rect 147404 567944 147456 567996
rect 157340 567944 157392 567996
rect 194784 567944 194836 567996
rect 302332 567944 302384 567996
rect 66352 567876 66404 567928
rect 121552 567876 121604 567928
rect 148784 567876 148836 567928
rect 161480 567876 161532 567928
rect 183652 567876 183704 567928
rect 301136 567876 301188 567928
rect 63500 567808 63552 567860
rect 123484 567808 123536 567860
rect 148876 567808 148928 567860
rect 164332 567808 164384 567860
rect 179420 567808 179472 567860
rect 300860 567808 300912 567860
rect 293960 567740 294012 567792
rect 319536 567740 319588 567792
rect 289820 567672 289872 567724
rect 314108 567672 314160 567724
rect 291200 567604 291252 567656
rect 314200 567604 314252 567656
rect 149796 567196 149848 567248
rect 151820 567196 151872 567248
rect 57060 566720 57112 566772
rect 62120 566720 62172 566772
rect 156604 566720 156656 566772
rect 213184 566720 213236 566772
rect 269120 566720 269172 566772
rect 317144 566720 317196 566772
rect 125692 566652 125744 566704
rect 211436 566652 211488 566704
rect 227720 566652 227772 566704
rect 300952 566652 301004 566704
rect 57520 566584 57572 566636
rect 82912 566584 82964 566636
rect 84200 566584 84252 566636
rect 122104 566584 122156 566636
rect 200120 566584 200172 566636
rect 302240 566584 302292 566636
rect 58532 566516 58584 566568
rect 110420 566516 110472 566568
rect 180984 566516 181036 566568
rect 301412 566516 301464 566568
rect 64880 566448 64932 566500
rect 122012 566448 122064 566500
rect 148508 566448 148560 566500
rect 160192 566448 160244 566500
rect 179512 566448 179564 566500
rect 301596 566448 301648 566500
rect 148692 565836 148744 565888
rect 150532 565836 150584 565888
rect 161572 565564 161624 565616
rect 178040 565564 178092 565616
rect 82728 565496 82780 565548
rect 89720 565496 89772 565548
rect 163044 565496 163096 565548
rect 183836 565496 183888 565548
rect 235448 565496 235500 565548
rect 248512 565496 248564 565548
rect 249064 565496 249116 565548
rect 271236 565496 271288 565548
rect 74632 565428 74684 565480
rect 96988 565428 97040 565480
rect 100208 565428 100260 565480
rect 115204 565428 115256 565480
rect 143540 565428 143592 565480
rect 166448 565428 166500 565480
rect 173900 565428 173952 565480
rect 189632 565428 189684 565480
rect 230480 565428 230532 565480
rect 259644 565428 259696 565480
rect 269764 565428 269816 565480
rect 282920 565428 282972 565480
rect 77024 565360 77076 565412
rect 84844 565360 84896 565412
rect 86040 565360 86092 565412
rect 108396 565360 108448 565412
rect 154672 565360 154724 565412
rect 181260 565360 181312 565412
rect 187792 565360 187844 565412
rect 198740 565360 198792 565412
rect 227812 565360 227864 565412
rect 265532 565360 265584 565412
rect 273352 565360 273404 565412
rect 296996 565360 297048 565412
rect 79876 565292 79928 565344
rect 114652 565292 114704 565344
rect 158720 565292 158772 565344
rect 192852 565292 192904 565344
rect 196624 565292 196676 565344
rect 210240 565292 210292 565344
rect 231952 565292 232004 565344
rect 279700 565292 279752 565344
rect 291844 565292 291896 565344
rect 300308 565292 300360 565344
rect 71320 565224 71372 565276
rect 109684 565224 109736 565276
rect 129740 565224 129792 565276
rect 163872 565224 163924 565276
rect 184204 565224 184256 565276
rect 213092 565224 213144 565276
rect 219440 565224 219492 565276
rect 268108 565224 268160 565276
rect 269212 565224 269264 565276
rect 307208 565224 307260 565276
rect 60280 565156 60332 565208
rect 104164 565156 104216 565208
rect 112444 565156 112496 565208
rect 117412 565156 117464 565208
rect 132592 565156 132644 565208
rect 187056 565156 187108 565208
rect 195244 565156 195296 565208
rect 212724 565156 212776 565208
rect 222292 565156 222344 565208
rect 273812 565156 273864 565208
rect 280160 565156 280212 565208
rect 322480 565156 322532 565208
rect 62856 565088 62908 565140
rect 108304 565088 108356 565140
rect 110512 565088 110564 565140
rect 120724 565088 120776 565140
rect 133972 565088 134024 565140
rect 207020 565088 207072 565140
rect 220820 565088 220872 565140
rect 239772 565088 239824 565140
rect 259460 565088 259512 565140
rect 321100 565088 321152 565140
rect 94504 564884 94556 564936
rect 102784 564884 102836 564936
rect 150348 564544 150400 564596
rect 151176 564544 151228 564596
rect 216680 564544 216732 564596
rect 220360 564544 220412 564596
rect 71780 564408 71832 564460
rect 73804 564408 73856 564460
rect 100760 564408 100812 564460
rect 102876 564408 102928 564460
rect 116584 564408 116636 564460
rect 120172 564408 120224 564460
rect 191104 564408 191156 564460
rect 195428 564408 195480 564460
rect 198004 564408 198056 564460
rect 201500 564408 201552 564460
rect 202144 564408 202196 564460
rect 204444 564408 204496 564460
rect 244924 564408 244976 564460
rect 250628 564408 250680 564460
rect 282184 564408 282236 564460
rect 288716 564408 288768 564460
rect 200212 563932 200264 563984
rect 239588 563932 239640 563984
rect 191840 563864 191892 563916
rect 238852 563864 238904 563916
rect 263600 563864 263652 563916
rect 322388 563864 322440 563916
rect 58900 563796 58952 563848
rect 91192 563796 91244 563848
rect 126980 563796 127032 563848
rect 211804 563796 211856 563848
rect 215392 563796 215444 563848
rect 301504 563796 301556 563848
rect 69020 563728 69072 563780
rect 123392 563728 123444 563780
rect 146852 563728 146904 563780
rect 165620 563728 165672 563780
rect 180892 563728 180944 563780
rect 301228 563728 301280 563780
rect 10324 563660 10376 563712
rect 321560 563660 321612 563712
rect 273260 562640 273312 562692
rect 322296 562640 322348 562692
rect 204260 562572 204312 562624
rect 239496 562572 239548 562624
rect 255320 562572 255372 562624
rect 324780 562572 324832 562624
rect 157524 562504 157576 562556
rect 212540 562504 212592 562556
rect 242900 562504 242952 562556
rect 318064 562504 318116 562556
rect 68744 562436 68796 562488
rect 106924 562436 106976 562488
rect 111892 562436 111944 562488
rect 123024 562436 123076 562488
rect 191932 562436 191984 562488
rect 273352 562436 273404 562488
rect 59452 562368 59504 562420
rect 75920 562368 75972 562420
rect 78772 562368 78824 562420
rect 121184 562368 121236 562420
rect 184940 562368 184992 562420
rect 294420 562368 294472 562420
rect 69112 562300 69164 562352
rect 114560 562300 114612 562352
rect 118700 562300 118752 562352
rect 154856 562300 154908 562352
rect 186320 562300 186372 562352
rect 302792 562300 302844 562352
rect 198740 561212 198792 561264
rect 239404 561212 239456 561264
rect 266452 561212 266504 561264
rect 307024 561212 307076 561264
rect 148232 561144 148284 561196
rect 158812 561144 158864 561196
rect 176660 561144 176712 561196
rect 217508 561144 217560 561196
rect 251180 561144 251232 561196
rect 323952 561144 324004 561196
rect 59268 561076 59320 561128
rect 92572 561076 92624 561128
rect 138020 561076 138072 561128
rect 211620 561076 211672 561128
rect 240140 561076 240192 561128
rect 313924 561076 313976 561128
rect 70400 561008 70452 561060
rect 121920 561008 121972 561060
rect 147036 561008 147088 561060
rect 168380 561008 168432 561060
rect 187700 561008 187752 561060
rect 301044 561008 301096 561060
rect 63592 560940 63644 560992
rect 122840 560940 122892 560992
rect 147312 560940 147364 560992
rect 175372 560940 175424 560992
rect 182180 560940 182232 560992
rect 301688 560940 301740 560992
rect 201500 559784 201552 559836
rect 256700 559784 256752 559836
rect 88432 559716 88484 559768
rect 103520 559716 103572 559768
rect 176752 559716 176804 559768
rect 244280 559716 244332 559768
rect 57244 559648 57296 559700
rect 89812 559648 89864 559700
rect 190460 559648 190512 559700
rect 277492 559648 277544 559700
rect 85672 559580 85724 559632
rect 121828 559580 121880 559632
rect 122840 559580 122892 559632
rect 211344 559580 211396 559632
rect 244280 559580 244332 559632
rect 319444 559580 319496 559632
rect 65064 559512 65116 559564
rect 123116 559512 123168 559564
rect 149060 559512 149112 559564
rect 160284 559512 160336 559564
rect 195980 559512 196032 559564
rect 302608 559512 302660 559564
rect 267740 558900 267792 558952
rect 321560 558900 321612 558952
rect 190552 558424 190604 558476
rect 222844 558424 222896 558476
rect 270500 558424 270552 558476
rect 309784 558424 309836 558476
rect 88432 558356 88484 558408
rect 104900 558356 104952 558408
rect 178040 558356 178092 558408
rect 236736 558356 236788 558408
rect 249800 558356 249852 558408
rect 307116 558356 307168 558408
rect 98644 558288 98696 558340
rect 123300 558288 123352 558340
rect 205640 558288 205692 558340
rect 285680 558288 285732 558340
rect 80060 558220 80112 558272
rect 120816 558220 120868 558272
rect 122932 558220 122984 558272
rect 211712 558220 211764 558272
rect 252560 558220 252612 558272
rect 323860 558220 323912 558272
rect 59544 558152 59596 558204
rect 100852 558152 100904 558204
rect 131120 558152 131172 558204
rect 187792 558152 187844 558204
rect 196072 558152 196124 558204
rect 302976 558152 303028 558204
rect 199200 557064 199252 557116
rect 232504 557064 232556 557116
rect 80980 556996 81032 557048
rect 121092 556996 121144 557048
rect 189908 556996 189960 557048
rect 238208 556996 238260 557048
rect 57428 556928 57480 556980
rect 81716 556928 81768 556980
rect 137192 556928 137244 556980
rect 212816 556928 212868 556980
rect 250812 556928 250864 556980
rect 323768 556928 323820 556980
rect 121092 556860 121144 556912
rect 198004 556860 198056 556912
rect 202236 556860 202288 556912
rect 302884 556860 302936 556912
rect 59084 556792 59136 556844
rect 102508 556792 102560 556844
rect 147220 556792 147272 556844
rect 174912 556792 174964 556844
rect 179144 556792 179196 556844
rect 291292 556792 291344 556844
rect 125600 555772 125652 555824
rect 126888 555772 126940 555824
rect 197820 555636 197872 555688
rect 216036 555636 216088 555688
rect 73160 555568 73212 555620
rect 107660 555568 107712 555620
rect 142620 555568 142672 555620
rect 213000 555568 213052 555620
rect 282368 555568 282420 555620
rect 305736 555568 305788 555620
rect 189172 555500 189224 555552
rect 282184 555500 282236 555552
rect 283748 555500 283800 555552
rect 312636 555500 312688 555552
rect 59176 555432 59228 555484
rect 108212 555432 108264 555484
rect 187056 555432 187108 555484
rect 302424 555432 302476 555484
rect 21364 554752 21416 554804
rect 321560 554752 321612 554804
rect 193496 554344 193548 554396
rect 217416 554344 217468 554396
rect 206376 554276 206428 554328
rect 262220 554276 262272 554328
rect 279516 554276 279568 554328
rect 311164 554276 311216 554328
rect 168380 554208 168432 554260
rect 210700 554208 210752 554260
rect 257988 554208 258040 554260
rect 321008 554208 321060 554260
rect 57796 554140 57848 554192
rect 103244 554140 103296 554192
rect 151176 554140 151228 554192
rect 163412 554140 163464 554192
rect 184940 554140 184992 554192
rect 235356 554140 235408 554192
rect 246488 554140 246540 554192
rect 312544 554140 312596 554192
rect 63132 554072 63184 554124
rect 110604 554072 110656 554124
rect 127624 554072 127676 554124
rect 202144 554072 202196 554124
rect 229284 554072 229336 554124
rect 303068 554072 303120 554124
rect 71688 554004 71740 554056
rect 121736 554004 121788 554056
rect 140504 554004 140556 554056
rect 196624 554004 196676 554056
rect 198556 554004 198608 554056
rect 291844 554004 291896 554056
rect 200212 553052 200264 553104
rect 201408 553052 201460 553104
rect 89812 552848 89864 552900
rect 91008 552848 91060 552900
rect 88432 552780 88484 552832
rect 89628 552780 89680 552832
rect 100760 552780 100812 552832
rect 101772 552780 101824 552832
rect 67640 552712 67692 552764
rect 68836 552712 68888 552764
rect 69020 552712 69072 552764
rect 70308 552712 70360 552764
rect 78680 552712 78732 552764
rect 79600 552712 79652 552764
rect 82452 552712 82504 552764
rect 76748 552644 76800 552696
rect 112444 552848 112496 552900
rect 116584 552712 116636 552764
rect 210792 552984 210844 553036
rect 213552 552984 213604 553036
rect 235264 552984 235316 553036
rect 173808 552916 173860 552968
rect 213368 552916 213420 552968
rect 260104 552916 260156 552968
rect 311256 552916 311308 552968
rect 122840 552712 122892 552764
rect 124036 552712 124088 552764
rect 124220 552712 124272 552764
rect 125416 552712 125468 552764
rect 126980 552712 127032 552764
rect 128268 552712 128320 552764
rect 211160 552848 211212 552900
rect 217876 552848 217928 552900
rect 269764 552848 269816 552900
rect 275192 552848 275244 552900
rect 316776 552848 316828 552900
rect 146300 552780 146352 552832
rect 213276 552780 213328 552832
rect 219440 552780 219492 552832
rect 220728 552780 220780 552832
rect 222200 552780 222252 552832
rect 222844 552780 222896 552832
rect 227720 552780 227772 552832
rect 228640 552780 228692 552832
rect 231860 552780 231912 552832
rect 232872 552780 232924 552832
rect 247960 552780 248012 552832
rect 324872 552780 324924 552832
rect 140780 552712 140832 552764
rect 141884 552712 141936 552764
rect 142160 552712 142212 552764
rect 143356 552712 143408 552764
rect 143540 552712 143592 552764
rect 144736 552712 144788 552764
rect 144920 552712 144972 552764
rect 146208 552712 146260 552764
rect 148508 552712 148560 552764
rect 172520 552712 172572 552764
rect 179420 552712 179472 552764
rect 180616 552712 180668 552764
rect 180892 552712 180944 552764
rect 181996 552712 182048 552764
rect 190460 552712 190512 552764
rect 191380 552712 191432 552764
rect 195980 552712 196032 552764
rect 197084 552712 197136 552764
rect 198740 552712 198792 552764
rect 199936 552712 199988 552764
rect 201500 552712 201552 552764
rect 202788 552712 202840 552764
rect 213920 552712 213972 552764
rect 215024 552712 215076 552764
rect 106280 552644 106332 552696
rect 107568 552644 107620 552696
rect 110420 552644 110472 552696
rect 111064 552644 111116 552696
rect 121828 552644 121880 552696
rect 129740 552644 129792 552696
rect 158720 552644 158772 552696
rect 159824 552644 159876 552696
rect 212172 552644 212224 552696
rect 302516 552712 302568 552764
rect 121460 552576 121512 552628
rect 122564 552576 122616 552628
rect 210700 552576 210752 552628
rect 301320 552644 301372 552696
rect 255320 552576 255372 552628
rect 256516 552576 256568 552628
rect 266360 552576 266412 552628
rect 267280 552576 267332 552628
rect 273260 552576 273312 552628
rect 274456 552576 274508 552628
rect 293960 552576 294012 552628
rect 295248 552576 295300 552628
rect 293132 552440 293184 552492
rect 316960 552440 317012 552492
rect 290924 552372 290976 552424
rect 316868 552372 316920 552424
rect 286692 552304 286744 552356
rect 313924 552304 313976 552356
rect 285220 552236 285272 552288
rect 317052 552236 317104 552288
rect 285956 552168 286008 552220
rect 319444 552168 319496 552220
rect 252928 552100 252980 552152
rect 322388 552100 322440 552152
rect 237932 552032 237984 552084
rect 322572 552032 322624 552084
rect 148416 551964 148468 552016
rect 149060 551964 149112 552016
rect 211436 551964 211488 552016
rect 214656 551964 214708 552016
rect 148600 551896 148652 551948
rect 149796 551896 149848 551948
rect 207112 551624 207164 551676
rect 220268 551624 220320 551676
rect 207848 551556 207900 551608
rect 229744 551556 229796 551608
rect 135444 551488 135496 551540
rect 144276 551488 144328 551540
rect 147680 551488 147732 551540
rect 191104 551488 191156 551540
rect 208584 551488 208636 551540
rect 238300 551488 238352 551540
rect 152648 551420 152700 551472
rect 211528 551420 211580 551472
rect 249432 551420 249484 551472
rect 301504 551420 301556 551472
rect 120448 551352 120500 551404
rect 130568 551352 130620 551404
rect 188528 551352 188580 551404
rect 253940 551352 253992 551404
rect 57612 551284 57664 551336
rect 77392 551284 77444 551336
rect 94596 551284 94648 551336
rect 123392 551284 123444 551336
rect 124680 551284 124732 551336
rect 210884 551284 210936 551336
rect 247224 551284 247276 551336
rect 301596 551284 301648 551336
rect 265900 551216 265952 551268
rect 307024 551216 307076 551268
rect 255872 551148 255924 551200
rect 304448 551148 304500 551200
rect 273076 551080 273128 551132
rect 321008 551080 321060 551132
rect 273720 551012 273772 551064
rect 323768 551012 323820 551064
rect 265164 550944 265216 550996
rect 318064 550944 318116 550996
rect 291660 550876 291712 550928
rect 316776 550876 316828 550928
rect 287336 550808 287388 550860
rect 317144 550808 317196 550860
rect 264428 550740 264480 550792
rect 322480 550740 322532 550792
rect 263048 550672 263100 550724
rect 322296 550672 322348 550724
rect 244372 550604 244424 550656
rect 324872 550604 324924 550656
rect 84844 550536 84896 550588
rect 86776 550536 86828 550588
rect 96068 550536 96120 550588
rect 98644 550536 98696 550588
rect 104164 550536 104216 550588
rect 105360 550536 105412 550588
rect 108304 550536 108356 550588
rect 109684 550536 109736 550588
rect 115204 550536 115256 550588
rect 116124 550536 116176 550588
rect 136180 550536 136232 550588
rect 140044 550536 140096 550588
rect 146944 550536 146996 550588
rect 148324 550536 148376 550588
rect 149888 550536 149940 550588
rect 151268 550536 151320 550588
rect 230020 550536 230072 550588
rect 231124 550536 231176 550588
rect 234344 550536 234396 550588
rect 236644 550536 236696 550588
rect 291200 550536 291252 550588
rect 292396 550536 292448 550588
rect 299572 550536 299624 550588
rect 304356 550536 304408 550588
rect 55128 550468 55180 550520
rect 67364 550468 67416 550520
rect 106924 550468 106976 550520
rect 108948 550468 109000 550520
rect 298836 550468 298888 550520
rect 304264 550468 304316 550520
rect 54944 550400 54996 550452
rect 88892 550400 88944 550452
rect 91100 550400 91152 550452
rect 96804 550400 96856 550452
rect 108396 550400 108448 550452
rect 111800 550400 111852 550452
rect 171324 550400 171376 550452
rect 173808 550400 173860 550452
rect 209228 550400 209280 550452
rect 217324 550400 217376 550452
rect 58716 550332 58768 550384
rect 95332 550332 95384 550384
rect 144092 550332 144144 550384
rect 146300 550332 146352 550384
rect 151084 550332 151136 550384
rect 153384 550332 153436 550384
rect 204260 550332 204312 550384
rect 215944 550332 215996 550384
rect 56508 550264 56560 550316
rect 83924 550264 83976 550316
rect 85304 550264 85356 550316
rect 121644 550264 121696 550316
rect 157800 550264 157852 550316
rect 167000 550264 167052 550316
rect 203524 550264 203576 550316
rect 220084 550264 220136 550316
rect 225052 550264 225104 550316
rect 235448 550264 235500 550316
rect 55036 550196 55088 550248
rect 93216 550196 93268 550248
rect 114008 550196 114060 550248
rect 125784 550196 125836 550248
rect 146116 550196 146168 550248
rect 156972 550196 157024 550248
rect 169852 550196 169904 550248
rect 175280 550196 175332 550248
rect 195612 550196 195664 550248
rect 214564 550196 214616 550248
rect 219992 550196 220044 550248
rect 233884 550196 233936 550248
rect 257252 550196 257304 550248
rect 300584 550196 300636 550248
rect 56416 550128 56468 550180
rect 98920 550128 98972 550180
rect 102784 550128 102836 550180
rect 106096 550128 106148 550180
rect 106832 550128 106884 550180
rect 124404 550128 124456 550180
rect 152004 550128 152056 550180
rect 167736 550128 167788 550180
rect 170588 550128 170640 550180
rect 195244 550128 195296 550180
rect 209964 550128 210016 550180
rect 228364 550128 228416 550180
rect 230756 550128 230808 550180
rect 244924 550128 244976 550180
rect 270868 550128 270920 550180
rect 322756 550128 322808 550180
rect 57704 550060 57756 550112
rect 99656 550060 99708 550112
rect 103980 550060 104032 550112
rect 124312 550060 124364 550112
rect 139032 550060 139084 550112
rect 184296 550060 184348 550112
rect 194232 550060 194284 550112
rect 220176 550060 220228 550112
rect 225788 550060 225840 550112
rect 241520 550060 241572 550112
rect 242256 550060 242308 550112
rect 323952 550060 324004 550112
rect 56324 549992 56376 550044
rect 73804 549992 73856 550044
rect 78128 549992 78180 550044
rect 122196 549992 122248 550044
rect 136916 549992 136968 550044
rect 156604 549992 156656 550044
rect 160100 549992 160152 550044
rect 172704 549992 172756 550044
rect 183468 549992 183520 550044
rect 231216 549992 231268 550044
rect 60372 549924 60424 549976
rect 116860 549924 116912 549976
rect 129004 549924 129056 549976
rect 137192 549924 137244 549976
rect 154120 549924 154172 549976
rect 204904 549924 204956 549976
rect 212816 549924 212868 549976
rect 249064 549924 249116 549976
rect 252284 549924 252336 549976
rect 293960 549924 294012 549976
rect 58624 549856 58676 549908
rect 117596 549856 117648 549908
rect 118976 549856 119028 549908
rect 128912 549856 128964 549908
rect 131856 549856 131908 549908
rect 144184 549856 144236 549908
rect 148968 549856 149020 549908
rect 171968 549856 172020 549908
rect 176292 549856 176344 549908
rect 238116 549856 238168 549908
rect 280160 549856 280212 549908
rect 301688 549856 301740 549908
rect 169760 549788 169812 549840
rect 173440 549788 173492 549840
rect 276572 549788 276624 549840
rect 300124 549788 300176 549840
rect 277308 549720 277360 549772
rect 300400 549720 300452 549772
rect 275928 549652 275980 549704
rect 302884 549652 302936 549704
rect 284484 549584 284536 549636
rect 319536 549584 319588 549636
rect 294512 549516 294564 549568
rect 319720 549516 319772 549568
rect 243636 549448 243688 549500
rect 287612 549448 287664 549500
rect 109776 549380 109828 549432
rect 114652 549380 114704 549432
rect 283104 549380 283156 549432
rect 295984 549448 296036 549500
rect 319628 549448 319680 549500
rect 322664 549380 322716 549432
rect 61660 549312 61712 549364
rect 64972 549312 65024 549364
rect 118240 549312 118292 549364
rect 124864 549312 124916 549364
rect 287888 549312 287940 549364
rect 300492 549312 300544 549364
rect 278044 549244 278096 549296
rect 300308 549244 300360 549296
rect 296720 548768 296772 548820
rect 319812 548768 319864 548820
rect 278780 548700 278832 548752
rect 300768 548700 300820 548752
rect 281632 548632 281684 548684
rect 287888 548632 287940 548684
rect 293960 548632 294012 548684
rect 321836 548632 321888 548684
rect 268752 548564 268804 548616
rect 300216 548564 300268 548616
rect 287612 548496 287664 548548
rect 322204 548496 322256 548548
rect 272340 548428 272392 548480
rect 304264 548428 304316 548480
rect 262312 548360 262364 548412
rect 324780 548360 324832 548412
rect 260840 548292 260892 548344
rect 323676 548292 323728 548344
rect 240048 548224 240100 548276
rect 302976 548224 303028 548276
rect 236460 548156 236512 548208
rect 302056 548156 302108 548208
rect 235816 548088 235868 548140
rect 254400 548088 254452 548140
rect 324688 548088 324740 548140
rect 323860 548020 323912 548072
rect 300768 542308 300820 542360
rect 321560 542308 321612 542360
rect 302608 539588 302660 539640
rect 320824 539588 320876 539640
rect 302056 536732 302108 536784
rect 321560 536732 321612 536784
rect 436744 527960 436796 528012
rect 436928 527960 436980 528012
rect 436376 527688 436428 527740
rect 436652 527688 436704 527740
rect 302976 527076 303028 527128
rect 321560 527076 321612 527128
rect 300492 522928 300544 522980
rect 436560 522928 436612 522980
rect 300400 522860 300452 522912
rect 436468 522860 436520 522912
rect 300584 522792 300636 522844
rect 436192 522792 436244 522844
rect 301780 522724 301832 522776
rect 436836 522724 436888 522776
rect 301872 522656 301924 522708
rect 433524 522656 433576 522708
rect 321100 522588 321152 522640
rect 436100 522588 436152 522640
rect 322756 522520 322808 522572
rect 436652 522520 436704 522572
rect 323952 522452 324004 522504
rect 436744 522452 436796 522504
rect 324872 522384 324924 522436
rect 325148 522384 325200 522436
rect 323584 521568 323636 521620
rect 342720 521568 342772 521620
rect 319444 521500 319496 521552
rect 495440 521500 495492 521552
rect 319812 521432 319864 521484
rect 459560 521432 459612 521484
rect 319628 521364 319680 521416
rect 457444 521364 457496 521416
rect 300308 521296 300360 521348
rect 436928 521296 436980 521348
rect 301688 521228 301740 521280
rect 436284 521228 436336 521280
rect 300124 521160 300176 521212
rect 420000 521160 420052 521212
rect 319536 521092 319588 521144
rect 433432 521092 433484 521144
rect 322388 521024 322440 521076
rect 433708 521024 433760 521076
rect 322572 520956 322624 521008
rect 433616 520956 433668 521008
rect 322664 520888 322716 520940
rect 433340 520888 433392 520940
rect 305644 520820 305696 520872
rect 374276 520820 374328 520872
rect 302884 520752 302936 520804
rect 356244 520752 356296 520804
rect 319720 520684 319772 520736
rect 500960 520684 501012 520736
rect 323676 520276 323728 520328
rect 318064 520208 318116 520260
rect 324688 520208 324740 520260
rect 347228 520208 347280 520260
rect 323860 520140 323912 520192
rect 338212 520140 338264 520192
rect 324596 520072 324648 520124
rect 334072 520072 334124 520124
rect 300216 520004 300268 520056
rect 393320 520004 393372 520056
rect 322296 519936 322348 519988
rect 406476 519936 406528 519988
rect 307024 519868 307076 519920
rect 388444 519868 388496 519920
rect 323768 519800 323820 519852
rect 401968 519800 402020 519852
rect 301596 519732 301648 519784
rect 365260 519732 365312 519784
rect 322480 519664 322532 519716
rect 379520 519664 379572 519716
rect 321008 519596 321060 519648
rect 369860 519596 369912 519648
rect 324504 519528 324556 519580
rect 351920 519528 351972 519580
rect 304264 519460 304316 519512
rect 415492 519460 415544 519512
rect 304448 519392 304500 519444
rect 411352 519392 411404 519444
rect 325148 519324 325200 519376
rect 424508 519324 424560 519376
rect 317144 518848 317196 518900
rect 476120 518848 476172 518900
rect 317052 518780 317104 518832
rect 470600 518780 470652 518832
rect 316776 518712 316828 518764
rect 457628 518712 457680 518764
rect 302976 518168 303028 518220
rect 576124 518168 576176 518220
rect 52368 517488 52420 517540
rect 57888 517488 57940 517540
rect 313924 517420 313976 517472
rect 512184 517420 512236 517472
rect 316960 517352 317012 517404
rect 512276 517352 512328 517404
rect 316868 517284 316920 517336
rect 488540 517284 488592 517336
rect 317236 517216 317288 517268
rect 465080 517216 465132 517268
rect 3424 514768 3476 514820
rect 11704 514768 11756 514820
rect 560944 511912 560996 511964
rect 580172 511912 580224 511964
rect 302240 495456 302292 495508
rect 520924 495456 520976 495508
rect 320824 489132 320876 489184
rect 580264 489132 580316 489184
rect 11704 488044 11756 488096
rect 360200 488044 360252 488096
rect 293976 487772 294028 487824
rect 294144 487772 294196 487824
rect 205824 487024 205876 487076
rect 206100 487024 206152 487076
rect 109500 486616 109552 486668
rect 204260 486616 204312 486668
rect 109408 486548 109460 486600
rect 205640 486548 205692 486600
rect 51908 486480 51960 486532
rect 99380 486480 99432 486532
rect 140872 486480 140924 486532
rect 199108 486480 199160 486532
rect 203616 486480 203668 486532
rect 356612 486480 356664 486532
rect 15844 486412 15896 486464
rect 383660 486412 383712 486464
rect 56416 485732 56468 485784
rect 81716 485732 81768 485784
rect 151268 485732 151320 485784
rect 211160 485732 211212 485784
rect 73896 485664 73948 485716
rect 102876 485664 102928 485716
rect 153936 485664 153988 485716
rect 212540 485664 212592 485716
rect 59912 485596 59964 485648
rect 91836 485596 91888 485648
rect 166172 485596 166224 485648
rect 211160 485596 211212 485648
rect 56508 485528 56560 485580
rect 89168 485528 89220 485580
rect 150440 485528 150492 485580
rect 69664 485460 69716 485512
rect 92296 485460 92348 485512
rect 152188 485460 152240 485512
rect 201408 485528 201460 485580
rect 211620 485528 211672 485580
rect 242072 485528 242124 485580
rect 356704 485528 356756 485580
rect 56324 485392 56376 485444
rect 88340 485392 88392 485444
rect 149428 485392 149480 485444
rect 191196 485392 191248 485444
rect 206192 485460 206244 485512
rect 240048 485460 240100 485512
rect 358268 485460 358320 485512
rect 204444 485392 204496 485444
rect 208308 485392 208360 485444
rect 217416 485392 217468 485444
rect 239680 485392 239732 485444
rect 358360 485392 358412 485444
rect 64144 485324 64196 485376
rect 72424 485324 72476 485376
rect 73896 485324 73948 485376
rect 106372 485324 106424 485376
rect 186320 485324 186372 485376
rect 193864 485324 193916 485376
rect 208952 485324 209004 485376
rect 218152 485324 218204 485376
rect 234528 485324 234580 485376
rect 363604 485324 363656 485376
rect 54668 485256 54720 485308
rect 102416 485256 102468 485308
rect 148232 485256 148284 485308
rect 51816 485188 51868 485240
rect 99748 485188 99800 485240
rect 139216 485188 139268 485240
rect 186320 485188 186372 485240
rect 195244 485256 195296 485308
rect 199384 485256 199436 485308
rect 197360 485188 197412 485240
rect 199844 485188 199896 485240
rect 217416 485256 217468 485308
rect 233240 485256 233292 485308
rect 366456 485256 366508 485308
rect 45468 485120 45520 485172
rect 105544 485120 105596 485172
rect 110328 485120 110380 485172
rect 164884 485120 164936 485172
rect 166264 485120 166316 485172
rect 202236 485120 202288 485172
rect 205456 485120 205508 485172
rect 219164 485188 219216 485240
rect 225604 485188 225656 485240
rect 358176 485188 358228 485240
rect 219072 485120 219124 485172
rect 219716 485120 219768 485172
rect 224040 485120 224092 485172
rect 360844 485120 360896 485172
rect 56232 485052 56284 485104
rect 90548 485052 90600 485104
rect 95424 485052 95476 485104
rect 167828 485052 167880 485104
rect 182272 485052 182324 485104
rect 208400 485052 208452 485104
rect 209504 485052 209556 485104
rect 221740 485052 221792 485104
rect 223488 485052 223540 485104
rect 371884 485052 371936 485104
rect 58624 484984 58676 485036
rect 81256 484984 81308 485036
rect 149888 484984 149940 485036
rect 197360 484984 197412 485036
rect 202696 484984 202748 485036
rect 210148 484984 210200 485036
rect 53656 484916 53708 484968
rect 74448 484916 74500 484968
rect 156604 484916 156656 484968
rect 166172 484916 166224 484968
rect 166264 484916 166316 484968
rect 201500 484916 201552 484968
rect 209044 484916 209096 484968
rect 219164 484916 219216 484968
rect 59176 484848 59228 484900
rect 69664 484848 69716 484900
rect 53288 484780 53340 484832
rect 68284 484712 68336 484764
rect 84384 484848 84436 484900
rect 139400 484848 139452 484900
rect 185584 484848 185636 484900
rect 191196 484848 191248 484900
rect 200488 484848 200540 484900
rect 157432 484780 157484 484832
rect 208400 484780 208452 484832
rect 155592 484712 155644 484764
rect 166264 484712 166316 484764
rect 167828 484712 167880 484764
rect 182824 484712 182876 484764
rect 77760 484644 77812 484696
rect 195152 484372 195204 484424
rect 197084 484372 197136 484424
rect 213368 484372 213420 484424
rect 214932 484372 214984 484424
rect 219992 484372 220044 484424
rect 222660 484372 222712 484424
rect 203708 484304 203760 484356
rect 209596 484304 209648 484356
rect 161572 484236 161624 484288
rect 162768 484236 162820 484288
rect 226616 484236 226668 484288
rect 227628 484236 227680 484288
rect 92572 484168 92624 484220
rect 93308 484168 93360 484220
rect 103520 484168 103572 484220
rect 104348 484168 104400 484220
rect 129832 484168 129884 484220
rect 130660 484168 130712 484220
rect 143632 484168 143684 484220
rect 143908 484168 143960 484220
rect 161480 484168 161532 484220
rect 161940 484168 161992 484220
rect 219532 484168 219584 484220
rect 219900 484168 219952 484220
rect 265164 484168 265216 484220
rect 265900 484168 265952 484220
rect 266452 484168 266504 484220
rect 267188 484168 267240 484220
rect 60740 484100 60792 484152
rect 61108 484100 61160 484152
rect 62120 484100 62172 484152
rect 62948 484100 63000 484152
rect 64880 484100 64932 484152
rect 65524 484100 65576 484152
rect 67732 484100 67784 484152
rect 68192 484100 68244 484152
rect 69020 484100 69072 484152
rect 69572 484100 69624 484152
rect 92480 484100 92532 484152
rect 92940 484100 92992 484152
rect 93860 484100 93912 484152
rect 94596 484100 94648 484152
rect 99472 484100 99524 484152
rect 100300 484100 100352 484152
rect 103612 484100 103664 484152
rect 103796 484100 103848 484152
rect 107660 484100 107712 484152
rect 107844 484100 107896 484152
rect 122840 484100 122892 484152
rect 123668 484100 123720 484152
rect 124312 484100 124364 484152
rect 124956 484100 125008 484152
rect 125600 484100 125652 484152
rect 126336 484100 126388 484152
rect 129924 484100 129976 484152
rect 130292 484100 130344 484152
rect 131120 484100 131172 484152
rect 132132 484100 132184 484152
rect 133880 484100 133932 484152
rect 134340 484100 134392 484152
rect 139400 484100 139452 484152
rect 140044 484100 140096 484152
rect 140872 484100 140924 484152
rect 141700 484100 141752 484152
rect 142160 484100 142212 484152
rect 142620 484100 142672 484152
rect 143540 484100 143592 484152
rect 144460 484100 144512 484152
rect 147680 484100 147732 484152
rect 148324 484100 148376 484152
rect 160100 484100 160152 484152
rect 160652 484100 160704 484152
rect 161572 484100 161624 484152
rect 162492 484100 162544 484152
rect 162860 484100 162912 484152
rect 163780 484100 163832 484152
rect 196716 484100 196768 484152
rect 196900 484100 196952 484152
rect 197452 484100 197504 484152
rect 198372 484100 198424 484152
rect 198740 484100 198792 484152
rect 198924 484100 198976 484152
rect 204444 484100 204496 484152
rect 205180 484100 205232 484152
rect 215392 484100 215444 484152
rect 216220 484100 216272 484152
rect 216772 484100 216824 484152
rect 217508 484100 217560 484152
rect 219624 484100 219676 484152
rect 220084 484100 220136 484152
rect 227720 484100 227772 484152
rect 228548 484100 228600 484152
rect 229100 484100 229152 484152
rect 229468 484100 229520 484152
rect 236000 484100 236052 484152
rect 236828 484100 236880 484152
rect 241520 484100 241572 484152
rect 242164 484100 242216 484152
rect 265072 484100 265124 484152
rect 265532 484100 265584 484152
rect 266360 484100 266412 484152
rect 266820 484100 266872 484152
rect 284300 484100 284352 484152
rect 284852 484100 284904 484152
rect 287060 484100 287112 484152
rect 287980 484100 288032 484152
rect 289912 484100 289964 484152
rect 290556 484100 290608 484152
rect 291292 484100 291344 484152
rect 291936 484100 291988 484152
rect 264980 484032 265032 484084
rect 265348 484032 265400 484084
rect 281448 484032 281500 484084
rect 60832 483964 60884 484016
rect 61660 483964 61712 484016
rect 286968 484032 287020 484084
rect 356888 484032 356940 484084
rect 376392 483964 376444 484016
rect 269028 483896 269080 483948
rect 370412 483896 370464 483948
rect 268016 483828 268068 483880
rect 377312 483828 377364 483880
rect 177304 483760 177356 483812
rect 205180 483760 205232 483812
rect 246028 483760 246080 483812
rect 369216 483760 369268 483812
rect 60648 483692 60700 483744
rect 80704 483692 80756 483744
rect 162768 483692 162820 483744
rect 215944 483692 215996 483744
rect 227904 483692 227956 483744
rect 362224 483692 362276 483744
rect 56784 483624 56836 483676
rect 113456 483624 113508 483676
rect 160008 483624 160060 483676
rect 214564 483624 214616 483676
rect 227628 483624 227680 483676
rect 370504 483624 370556 483676
rect 201500 483488 201552 483540
rect 201684 483488 201736 483540
rect 223580 483352 223632 483404
rect 224132 483352 224184 483404
rect 50436 482944 50488 482996
rect 97172 482944 97224 482996
rect 50528 482876 50580 482928
rect 98460 482876 98512 482928
rect 299388 482876 299440 482928
rect 364064 482876 364116 482928
rect 48044 482808 48096 482860
rect 98000 482808 98052 482860
rect 284760 482808 284812 482860
rect 359832 482808 359884 482860
rect 48136 482740 48188 482792
rect 111708 482740 111760 482792
rect 177120 482740 177172 482792
rect 203616 482740 203668 482792
rect 280068 482740 280120 482792
rect 361304 482740 361356 482792
rect 46664 482672 46716 482724
rect 111248 482672 111300 482724
rect 173440 482672 173492 482724
rect 216036 482672 216088 482724
rect 278688 482672 278740 482724
rect 362684 482672 362736 482724
rect 50620 482604 50672 482656
rect 115664 482604 115716 482656
rect 138480 482604 138532 482656
rect 46388 482536 46440 482588
rect 112076 482536 112128 482588
rect 140780 482536 140832 482588
rect 141332 482536 141384 482588
rect 165528 482604 165580 482656
rect 214656 482604 214708 482656
rect 272432 482604 272484 482656
rect 369676 482604 369728 482656
rect 197176 482536 197228 482588
rect 242900 482536 242952 482588
rect 243084 482536 243136 482588
rect 257528 482536 257580 482588
rect 362500 482536 362552 482588
rect 49056 482468 49108 482520
rect 115204 482468 115256 482520
rect 135720 482468 135772 482520
rect 197912 482468 197964 482520
rect 261392 482468 261444 482520
rect 369492 482468 369544 482520
rect 46296 482400 46348 482452
rect 112536 482400 112588 482452
rect 138848 482400 138900 482452
rect 201776 482400 201828 482452
rect 255228 482400 255280 482452
rect 369584 482400 369636 482452
rect 46756 482332 46808 482384
rect 119620 482332 119672 482384
rect 137928 482332 137980 482384
rect 203156 482332 203208 482384
rect 244648 482332 244700 482384
rect 372068 482332 372120 482384
rect 57244 482264 57296 482316
rect 135904 482264 135956 482316
rect 137560 482264 137612 482316
rect 204628 482264 204680 482316
rect 248328 482264 248380 482316
rect 378784 482264 378836 482316
rect 51632 482196 51684 482248
rect 97540 482196 97592 482248
rect 54576 482128 54628 482180
rect 96712 482128 96764 482180
rect 58808 482060 58860 482112
rect 96252 482060 96304 482112
rect 125692 481992 125744 482044
rect 125876 481992 125928 482044
rect 289728 481312 289780 481364
rect 372436 481312 372488 481364
rect 270040 481244 270092 481296
rect 358636 481244 358688 481296
rect 262220 481176 262272 481228
rect 262588 481176 262640 481228
rect 270408 481176 270460 481228
rect 359464 481176 359516 481228
rect 189172 481108 189224 481160
rect 189356 481108 189408 481160
rect 251364 481108 251416 481160
rect 251548 481108 251600 481160
rect 271788 481108 271840 481160
rect 377220 481108 377272 481160
rect 74724 481040 74776 481092
rect 74908 481040 74960 481092
rect 168564 481040 168616 481092
rect 168748 481040 168800 481092
rect 176016 481040 176068 481092
rect 209228 481040 209280 481092
rect 212724 481040 212776 481092
rect 212908 481040 212960 481092
rect 244096 481040 244148 481092
rect 363696 481040 363748 481092
rect 57796 480972 57848 481024
rect 114284 480972 114336 481024
rect 160560 480972 160612 481024
rect 211804 480972 211856 481024
rect 253112 480972 253164 481024
rect 374828 480972 374880 481024
rect 3700 480904 3752 480956
rect 434904 480904 434956 480956
rect 70400 480836 70452 480888
rect 70860 480836 70912 480888
rect 74632 480836 74684 480888
rect 75276 480836 75328 480888
rect 75920 480836 75972 480888
rect 76564 480836 76616 480888
rect 81532 480836 81584 480888
rect 82268 480836 82320 480888
rect 82912 480836 82964 480888
rect 83556 480836 83608 480888
rect 84292 480836 84344 480888
rect 84936 480836 84988 480888
rect 86960 480836 87012 480888
rect 87604 480836 87656 480888
rect 88432 480836 88484 480888
rect 89260 480836 89312 480888
rect 167092 480836 167144 480888
rect 167736 480836 167788 480888
rect 168380 480836 168432 480888
rect 169116 480836 169168 480888
rect 169760 480836 169812 480888
rect 170036 480836 170088 480888
rect 173900 480836 173952 480888
rect 174268 480836 174320 480888
rect 179420 480836 179472 480888
rect 180064 480836 180116 480888
rect 182272 480836 182324 480888
rect 183100 480836 183152 480888
rect 186320 480836 186372 480888
rect 187148 480836 187200 480888
rect 205824 480836 205876 480888
rect 206468 480836 206520 480888
rect 207204 480836 207256 480888
rect 207572 480836 207624 480888
rect 209780 480836 209832 480888
rect 209964 480836 210016 480888
rect 212540 480836 212592 480888
rect 213460 480836 213512 480888
rect 248420 480836 248472 480888
rect 249156 480836 249208 480888
rect 249892 480836 249944 480888
rect 250076 480836 250128 480888
rect 251180 480836 251232 480888
rect 251916 480836 251968 480888
rect 253940 480836 253992 480888
rect 254124 480836 254176 480888
rect 262312 480836 262364 480888
rect 262864 480836 262916 480888
rect 292580 480836 292632 480888
rect 293316 480836 293368 480888
rect 293960 480836 294012 480888
rect 294604 480836 294656 480888
rect 295524 480836 295576 480888
rect 296260 480836 296312 480888
rect 70492 480768 70544 480820
rect 71228 480768 71280 480820
rect 131212 480632 131264 480684
rect 131580 480632 131632 480684
rect 171140 480292 171192 480344
rect 171692 480292 171744 480344
rect 51724 480156 51776 480208
rect 116124 480156 116176 480208
rect 292764 480156 292816 480208
rect 368296 480156 368348 480208
rect 47400 480088 47452 480140
rect 117596 480088 117648 480140
rect 281724 480088 281776 480140
rect 359648 480088 359700 480140
rect 59636 480020 59688 480072
rect 129924 480020 129976 480072
rect 297732 480020 297784 480072
rect 376576 480020 376628 480072
rect 48964 479952 49016 480004
rect 121552 479952 121604 480004
rect 278872 479952 278924 480004
rect 364156 479952 364208 480004
rect 49148 479884 49200 479936
rect 127716 479884 127768 479936
rect 275192 479884 275244 479936
rect 370320 479884 370372 479936
rect 42524 479816 42576 479868
rect 122932 479816 122984 479868
rect 260932 479816 260984 479868
rect 368020 479816 368072 479868
rect 42432 479748 42484 479800
rect 123300 479748 123352 479800
rect 265256 479748 265308 479800
rect 373448 479748 373500 479800
rect 48872 479680 48924 479732
rect 129740 479680 129792 479732
rect 254492 479680 254544 479732
rect 366732 479680 366784 479732
rect 42340 479612 42392 479664
rect 124588 479612 124640 479664
rect 253204 479612 253256 479664
rect 374920 479612 374972 479664
rect 46112 479544 46164 479596
rect 129004 479544 129056 479596
rect 158996 479544 159048 479596
rect 207664 479544 207716 479596
rect 242992 479544 243044 479596
rect 366548 479544 366600 479596
rect 62396 479476 62448 479528
rect 199200 479476 199252 479528
rect 246488 479476 246540 479528
rect 369308 479476 369360 479528
rect 54484 479408 54536 479460
rect 117412 479408 117464 479460
rect 53288 479340 53340 479392
rect 116216 479340 116268 479392
rect 53380 479272 53432 479324
rect 116676 479272 116728 479324
rect 85580 479136 85632 479188
rect 86316 479136 86368 479188
rect 169852 478728 169904 478780
rect 170404 478728 170456 478780
rect 291476 478592 291528 478644
rect 361396 478592 361448 478644
rect 288900 478524 288952 478576
rect 361488 478524 361540 478576
rect 298468 478456 298520 478508
rect 379244 478456 379296 478508
rect 178132 478252 178184 478304
rect 210700 478252 210752 478304
rect 238208 478252 238260 478304
rect 247408 478320 247460 478372
rect 160192 478184 160244 478236
rect 203524 478184 203576 478236
rect 249800 478184 249852 478236
rect 250536 478184 250588 478236
rect 275652 478388 275704 478440
rect 373724 478388 373776 478440
rect 260196 478320 260248 478372
rect 370780 478320 370832 478372
rect 365076 478252 365128 478304
rect 376024 478184 376076 478236
rect 85672 478116 85724 478168
rect 85856 478116 85908 478168
rect 146300 478116 146352 478168
rect 218704 478116 218756 478168
rect 238760 478116 238812 478168
rect 378876 478116 378928 478168
rect 273352 477844 273404 477896
rect 273812 477844 273864 477896
rect 277400 477844 277452 477896
rect 277860 477844 277912 477896
rect 78772 477640 78824 477692
rect 79140 477640 79192 477692
rect 59728 477436 59780 477488
rect 133880 477436 133932 477488
rect 46848 477368 46900 477420
rect 122840 477368 122892 477420
rect 207112 477368 207164 477420
rect 207756 477368 207808 477420
rect 291292 477368 291344 477420
rect 365536 477368 365588 477420
rect 57336 477300 57388 477352
rect 135996 477300 136048 477352
rect 276572 477300 276624 477352
rect 358728 477300 358780 477352
rect 55772 477232 55824 477284
rect 134708 477232 134760 477284
rect 274732 477232 274784 477284
rect 365444 477232 365496 477284
rect 50160 477164 50212 477216
rect 131304 477164 131356 477216
rect 264244 477164 264296 477216
rect 362592 477164 362644 477216
rect 47860 477096 47912 477148
rect 129832 477096 129884 477148
rect 263600 477096 263652 477148
rect 363972 477096 364024 477148
rect 48780 477028 48832 477080
rect 133420 477028 133472 477080
rect 263692 477028 263744 477080
rect 365352 477028 365404 477080
rect 46204 476960 46256 477012
rect 132592 476960 132644 477012
rect 204536 476960 204588 477012
rect 217324 476960 217376 477012
rect 259736 476960 259788 477012
rect 363880 476960 363932 477012
rect 43996 476892 44048 476944
rect 132500 476892 132552 476944
rect 188068 476892 188120 476944
rect 207756 476892 207808 476944
rect 258540 476892 258592 476944
rect 368112 476892 368164 476944
rect 45008 476824 45060 476876
rect 133972 476824 134024 476876
rect 185768 476824 185820 476876
rect 213276 476824 213328 476876
rect 246120 476824 246172 476876
rect 362408 476824 362460 476876
rect 44732 476756 44784 476808
rect 143724 476756 143776 476808
rect 164608 476756 164660 476808
rect 211896 476756 211948 476808
rect 244464 476756 244516 476808
rect 373264 476756 373316 476808
rect 57152 476688 57204 476740
rect 131212 476688 131264 476740
rect 58440 476620 58492 476672
rect 131120 476620 131172 476672
rect 58532 476552 58584 476604
rect 128452 476552 128504 476604
rect 175280 476416 175332 476468
rect 176108 476416 176160 476468
rect 278780 475804 278832 475856
rect 357072 475804 357124 475856
rect 270868 475736 270920 475788
rect 364248 475736 364300 475788
rect 274640 475668 274692 475720
rect 368388 475668 368440 475720
rect 187792 475600 187844 475652
rect 200948 475600 201000 475652
rect 259460 475600 259512 475652
rect 372252 475600 372304 475652
rect 179604 475532 179656 475584
rect 219072 475532 219124 475584
rect 236460 475532 236512 475584
rect 362316 475532 362368 475584
rect 162952 475464 163004 475516
rect 206376 475464 206428 475516
rect 232412 475464 232464 475516
rect 367744 475464 367796 475516
rect 168656 475396 168708 475448
rect 213184 475396 213236 475448
rect 237472 475396 237524 475448
rect 376116 475396 376168 475448
rect 61016 475328 61068 475380
rect 199568 475328 199620 475380
rect 206100 475328 206152 475380
rect 217692 475328 217744 475380
rect 229192 475328 229244 475380
rect 369124 475328 369176 475380
rect 45376 474512 45428 474564
rect 73896 474512 73948 474564
rect 54760 474444 54812 474496
rect 101588 474444 101640 474496
rect 289912 474444 289964 474496
rect 367008 474444 367060 474496
rect 53196 474376 53248 474428
rect 99932 474376 99984 474428
rect 290188 474376 290240 474428
rect 374460 474376 374512 474428
rect 57428 474308 57480 474360
rect 103704 474308 103756 474360
rect 178040 474308 178092 474360
rect 202144 474308 202196 474360
rect 273444 474308 273496 474360
rect 360752 474308 360804 474360
rect 50344 474240 50396 474292
rect 98644 474240 98696 474292
rect 172060 474240 172112 474292
rect 210516 474240 210568 474292
rect 257620 474240 257672 474292
rect 366824 474240 366876 474292
rect 51540 474172 51592 474224
rect 99472 474172 99524 474224
rect 158720 474172 158772 474224
rect 209044 474172 209096 474224
rect 262404 474172 262456 474224
rect 373540 474172 373592 474224
rect 57704 474104 57756 474156
rect 113548 474104 113600 474156
rect 153200 474104 153252 474156
rect 218796 474104 218848 474156
rect 244372 474104 244424 474156
rect 360936 474104 360988 474156
rect 45284 474036 45336 474088
rect 106372 474036 106424 474088
rect 139492 474036 139544 474088
rect 207296 474036 207348 474088
rect 240140 474036 240192 474088
rect 369400 474036 369452 474088
rect 59360 473968 59412 474020
rect 180156 473968 180208 474020
rect 186412 473968 186464 474020
rect 212080 473968 212132 474020
rect 240784 473968 240836 474020
rect 374644 473968 374696 474020
rect 291200 473152 291252 473204
rect 357164 473152 357216 473204
rect 280160 473084 280212 473136
rect 366272 473084 366324 473136
rect 273352 473016 273404 473068
rect 362868 473016 362920 473068
rect 262312 472948 262364 473000
rect 372344 472948 372396 473000
rect 258172 472880 258224 472932
rect 370872 472880 370924 472932
rect 58716 472812 58768 472864
rect 110604 472812 110656 472864
rect 241612 472812 241664 472864
rect 376208 472812 376260 472864
rect 45192 472744 45244 472796
rect 105636 472744 105688 472796
rect 226340 472744 226392 472796
rect 364984 472744 365036 472796
rect 45100 472676 45152 472728
rect 104992 472676 105044 472728
rect 175372 472676 175424 472728
rect 210792 472676 210844 472728
rect 237380 472676 237432 472728
rect 378968 472676 379020 472728
rect 43444 472608 43496 472660
rect 103612 472608 103664 472660
rect 179512 472608 179564 472660
rect 216220 472608 216272 472660
rect 227260 472608 227312 472660
rect 371976 472608 372028 472660
rect 50896 471928 50948 471980
rect 81900 471928 81952 471980
rect 185032 471928 185084 471980
rect 206560 471928 206612 471980
rect 295892 471928 295944 471980
rect 369768 471928 369820 471980
rect 53564 471860 53616 471912
rect 84476 471860 84528 471912
rect 189724 471860 189776 471912
rect 215024 471860 215076 471912
rect 295524 471860 295576 471912
rect 370228 471860 370280 471912
rect 50804 471792 50856 471844
rect 82820 471792 82872 471844
rect 191012 471792 191064 471844
rect 217416 471792 217468 471844
rect 295432 471792 295484 471844
rect 371240 471792 371292 471844
rect 51448 471724 51500 471776
rect 84292 471724 84344 471776
rect 181444 471724 181496 471776
rect 209320 471724 209372 471776
rect 288440 471724 288492 471776
rect 364892 471724 364944 471776
rect 53656 471656 53708 471708
rect 85764 471656 85816 471708
rect 182732 471656 182784 471708
rect 210884 471656 210936 471708
rect 296720 471656 296772 471708
rect 373816 471656 373868 471708
rect 50712 471588 50764 471640
rect 82912 471588 82964 471640
rect 182272 471588 182324 471640
rect 216312 471588 216364 471640
rect 298100 471588 298152 471640
rect 375380 471588 375432 471640
rect 49424 471520 49476 471572
rect 83188 471520 83240 471572
rect 161664 471520 161716 471572
rect 210608 471520 210660 471572
rect 295340 471520 295392 471572
rect 377128 471520 377180 471572
rect 58900 471452 58952 471504
rect 95516 471452 95568 471504
rect 140964 471452 141016 471504
rect 200396 471452 200448 471504
rect 286140 471452 286192 471504
rect 377956 471452 378008 471504
rect 53104 471384 53156 471436
rect 100760 471384 100812 471436
rect 140872 471384 140924 471436
rect 195244 471384 195296 471436
rect 195336 471384 195388 471436
rect 200488 471384 200540 471436
rect 287152 471384 287204 471436
rect 379336 471384 379388 471436
rect 57520 471316 57572 471368
rect 114744 471316 114796 471368
rect 124220 471316 124272 471368
rect 196900 471316 196952 471368
rect 255412 471316 255464 471368
rect 358452 471316 358504 471368
rect 53012 471248 53064 471300
rect 100852 471248 100904 471300
rect 108212 471248 108264 471300
rect 202880 471248 202932 471300
rect 251364 471248 251416 471300
rect 366640 471248 366692 471300
rect 44916 471180 44968 471232
rect 65064 471180 65116 471232
rect 182364 471180 182416 471232
rect 203708 471180 203760 471232
rect 287520 471180 287572 471232
rect 359556 471180 359608 471232
rect 44824 471112 44876 471164
rect 64880 471112 64932 471164
rect 185584 471112 185636 471164
rect 205916 471112 205968 471164
rect 299480 471112 299532 471164
rect 364800 471112 364852 471164
rect 47768 471044 47820 471096
rect 64972 471044 65024 471096
rect 195244 471044 195296 471096
rect 201868 471044 201920 471096
rect 193864 470976 193916 471028
rect 195336 470976 195388 471028
rect 289820 470500 289872 470552
rect 360660 470500 360712 470552
rect 283104 470432 283156 470484
rect 358084 470432 358136 470484
rect 282920 470364 282972 470416
rect 359924 470364 359976 470416
rect 283012 470296 283064 470348
rect 360016 470296 360068 470348
rect 287060 470228 287112 470280
rect 367560 470228 367612 470280
rect 285772 470160 285824 470212
rect 373908 470160 373960 470212
rect 281540 470092 281592 470144
rect 371148 470092 371200 470144
rect 270500 470024 270552 470076
rect 362776 470024 362828 470076
rect 284392 469956 284444 470008
rect 377496 469956 377548 470008
rect 172612 469888 172664 469940
rect 205088 469888 205140 469940
rect 284300 469888 284352 469940
rect 377588 469888 377640 469940
rect 57612 469820 57664 469872
rect 111984 469820 112036 469872
rect 160100 469820 160152 469872
rect 202328 469820 202380 469872
rect 281632 469820 281684 469872
rect 379888 469820 379940 469872
rect 51356 469140 51408 469192
rect 68284 469140 68336 469192
rect 192024 469140 192076 469192
rect 213092 469140 213144 469192
rect 266360 469140 266412 469192
rect 359740 469140 359792 469192
rect 49608 469072 49660 469124
rect 70584 469072 70636 469124
rect 193404 469072 193456 469124
rect 217600 469072 217652 469124
rect 271972 469072 272024 469124
rect 366180 469072 366232 469124
rect 54944 469004 54996 469056
rect 85672 469004 85724 469056
rect 175280 469004 175332 469056
rect 206652 469004 206704 469056
rect 266544 469004 266596 469056
rect 361212 469004 361264 469056
rect 56048 468936 56100 468988
rect 87144 468936 87196 468988
rect 180892 468936 180944 468988
rect 212356 468936 212408 468988
rect 265164 468936 265216 468988
rect 361120 468936 361172 468988
rect 55036 468868 55088 468920
rect 86960 468868 87012 468920
rect 179420 468868 179472 468920
rect 214748 468868 214800 468920
rect 276020 468868 276072 468920
rect 374368 468868 374420 468920
rect 54852 468800 54904 468852
rect 88524 468800 88576 468852
rect 167184 468800 167236 468852
rect 209136 468800 209188 468852
rect 267740 468800 267792 468852
rect 369032 468800 369084 468852
rect 52092 468732 52144 468784
rect 85580 468732 85632 468784
rect 142344 468732 142396 468784
rect 199016 468732 199068 468784
rect 255320 468732 255372 468784
rect 356796 468732 356848 468784
rect 53472 468664 53524 468716
rect 87052 468664 87104 468716
rect 139400 468664 139452 468716
rect 197268 468664 197320 468716
rect 254032 468664 254084 468716
rect 358544 468664 358596 468716
rect 49332 468596 49384 468648
rect 92572 468596 92624 468648
rect 109040 468596 109092 468648
rect 197728 468596 197780 468648
rect 266452 468596 266504 468648
rect 375288 468596 375340 468648
rect 49240 468528 49292 468580
rect 93952 468528 94004 468580
rect 107752 468528 107804 468580
rect 197636 468528 197688 468580
rect 249984 468528 250036 468580
rect 365168 468528 365220 468580
rect 43352 468460 43404 468512
rect 103520 468460 103572 468512
rect 107660 468460 107712 468512
rect 201684 468460 201736 468512
rect 249892 468460 249944 468512
rect 373356 468460 373408 468512
rect 47676 468392 47728 468444
rect 63592 468392 63644 468444
rect 191932 468392 191984 468444
rect 211620 468392 211672 468444
rect 294052 468392 294104 468444
rect 375748 468392 375800 468444
rect 192116 468324 192168 468376
rect 210056 468324 210108 468376
rect 186320 468256 186372 468308
rect 200856 468256 200908 468308
rect 80704 467780 80756 467832
rect 178040 467780 178092 467832
rect 292672 467576 292724 467628
rect 357992 467576 358044 467628
rect 277492 467508 277544 467560
rect 367652 467508 367704 467560
rect 189172 467440 189224 467492
rect 200764 467440 200816 467492
rect 273260 467440 273312 467492
rect 363512 467440 363564 467492
rect 189080 467372 189132 467424
rect 202512 467372 202564 467424
rect 256700 467372 256752 467424
rect 361028 467372 361080 467424
rect 44088 467304 44140 467356
rect 70492 467304 70544 467356
rect 184940 467304 184992 467356
rect 212172 467304 212224 467356
rect 251272 467304 251324 467356
rect 365260 467304 365312 467356
rect 42248 467236 42300 467288
rect 73804 467236 73856 467288
rect 180156 467236 180208 467288
rect 218060 467236 218112 467288
rect 260840 467236 260892 467288
rect 376300 467236 376352 467288
rect 41328 467168 41380 467220
rect 93860 467168 93912 467220
rect 164240 467168 164292 467220
rect 218888 467168 218940 467220
rect 258080 467168 258132 467220
rect 373632 467168 373684 467220
rect 47952 467100 48004 467152
rect 106464 467100 106516 467152
rect 151820 467100 151872 467152
rect 210424 467100 210476 467152
rect 251180 467100 251232 467152
rect 366916 467100 366968 467152
rect 339408 466556 339460 466608
rect 361580 466556 361632 466608
rect 498476 466556 498528 466608
rect 517888 466556 517940 466608
rect 178040 466488 178092 466540
rect 190920 466420 190972 466472
rect 207020 466420 207072 466472
rect 218060 466488 218112 466540
rect 218244 466488 218296 466540
rect 339776 466488 339828 466540
rect 356980 466488 357032 466540
rect 499764 466488 499816 466540
rect 212816 466420 212868 466472
rect 338488 466420 338540 466472
rect 339408 466420 339460 466472
rect 351000 466420 351052 466472
rect 362960 466420 363012 466472
rect 510896 466488 510948 466540
rect 517520 466488 517572 466540
rect 517796 466420 517848 466472
rect 52000 466352 52052 466404
rect 75920 466352 75972 466404
rect 182180 466352 182232 466404
rect 202420 466352 202472 466404
rect 213828 466352 213880 466404
rect 221004 466352 221056 466404
rect 264980 466352 265032 466404
rect 368204 466352 368256 466404
rect 55680 466284 55732 466336
rect 77484 466284 77536 466336
rect 187700 466284 187752 466336
rect 211528 466284 211580 466336
rect 269120 466284 269172 466336
rect 372528 466284 372580 466336
rect 191840 466216 191892 466268
rect 215852 466216 215904 466268
rect 262220 466216 262272 466268
rect 379060 466216 379112 466268
rect 54392 466148 54444 466200
rect 62120 466148 62172 466200
rect 180800 466148 180852 466200
rect 206744 466148 206796 466200
rect 249800 466148 249852 466200
rect 367928 466148 367980 466200
rect 59268 466080 59320 466132
rect 67640 466080 67692 466132
rect 173992 466080 174044 466132
rect 203800 466080 203852 466132
rect 248512 466080 248564 466132
rect 370688 466080 370740 466132
rect 54300 466012 54352 466064
rect 63500 466012 63552 466064
rect 176660 466012 176712 466064
rect 209412 466012 209464 466064
rect 248420 466012 248472 466064
rect 372160 466012 372212 466064
rect 43260 465944 43312 465996
rect 60832 465944 60884 465996
rect 164884 465944 164936 465996
rect 200304 465944 200356 465996
rect 253940 465944 253992 465996
rect 379152 465944 379204 465996
rect 52276 465876 52328 465928
rect 70400 465876 70452 465928
rect 173900 465876 173952 465928
rect 214840 465876 214892 465928
rect 241520 465876 241572 465928
rect 367836 465876 367888 465928
rect 42156 465808 42208 465860
rect 60740 465808 60792 465860
rect 140780 465808 140832 465860
rect 203248 465808 203300 465860
rect 244280 465808 244332 465860
rect 370596 465808 370648 465860
rect 51448 465740 51500 465792
rect 52184 465740 52236 465792
rect 53748 465740 53800 465792
rect 74724 465740 74776 465792
rect 142252 465740 142304 465792
rect 207388 465740 207440 465792
rect 236000 465740 236052 465792
rect 363788 465740 363840 465792
rect 42708 465672 42760 465724
rect 66352 465672 66404 465724
rect 72424 465672 72476 465724
rect 198924 465672 198976 465724
rect 209688 465672 209740 465724
rect 220912 465672 220964 465724
rect 242900 465672 242952 465724
rect 374736 465672 374788 465724
rect 190552 465604 190604 465656
rect 199476 465604 199528 465656
rect 194600 465536 194652 465588
rect 213000 465604 213052 465656
rect 277400 465604 277452 465656
rect 364708 465604 364760 465656
rect 285680 465536 285732 465588
rect 357900 465536 357952 465588
rect 193312 465468 193364 465520
rect 203892 465468 203944 465520
rect 198924 465060 198976 465112
rect 358820 465060 358872 465112
rect 518900 465060 518952 465112
rect 51356 464992 51408 465044
rect 52000 464992 52052 465044
rect 197176 464992 197228 465044
rect 200580 464992 200632 465044
rect 207480 464992 207532 465044
rect 207940 464992 207992 465044
rect 190460 464720 190512 464772
rect 208768 464720 208820 464772
rect 59084 464652 59136 464704
rect 89904 464652 89956 464704
rect 183652 464652 183704 464704
rect 205272 464652 205324 464704
rect 58992 464584 59044 464636
rect 92480 464584 92532 464636
rect 183560 464584 183612 464636
rect 207848 464584 207900 464636
rect 55864 464516 55916 464568
rect 102324 464516 102376 464568
rect 193220 464516 193272 464568
rect 217784 464516 217836 464568
rect 52920 464448 52972 464500
rect 121460 464448 121512 464500
rect 126980 464448 127032 464500
rect 197820 464448 197872 464500
rect 57060 464380 57112 464432
rect 128360 464380 128412 464432
rect 142160 464380 142212 464432
rect 198004 464380 198056 464432
rect 293960 464380 294012 464432
rect 375012 464380 375064 464432
rect 55956 464312 56008 464364
rect 130016 464312 130068 464364
rect 136640 464312 136692 464364
rect 199292 464312 199344 464364
rect 271880 464312 271932 464364
rect 371792 464312 371844 464364
rect 46020 464244 46072 464296
rect 207940 464244 207992 464296
rect 207940 422900 207992 422952
rect 217968 422900 218020 422952
rect 55680 418208 55732 418260
rect 57152 418208 57204 418260
rect 55772 418140 55824 418192
rect 56876 418140 56928 418192
rect 46020 418072 46072 418124
rect 56968 418072 57020 418124
rect 207204 417460 207256 417512
rect 216680 417460 216732 417512
rect 206836 417392 206888 417444
rect 219624 417392 219676 417444
rect 357900 417392 357952 417444
rect 376944 417392 376996 417444
rect 44640 416780 44692 416832
rect 57888 416780 57940 416832
rect 205824 416712 205876 416764
rect 207940 416712 207992 416764
rect 55680 415352 55732 415404
rect 57060 415352 57112 415404
rect 57152 415352 57204 415404
rect 58440 415352 58492 415404
rect 207940 414808 207992 414860
rect 217140 414808 217192 414860
rect 208124 414740 208176 414792
rect 216864 414740 216916 414792
rect 206928 414672 206980 414724
rect 216772 414672 216824 414724
rect 359832 414672 359884 414724
rect 377680 414672 377732 414724
rect 47584 413992 47636 414044
rect 57888 413992 57940 414044
rect 57244 413924 57296 413976
rect 58440 413924 58492 413976
rect 205732 413244 205784 413296
rect 216864 413244 216916 413296
rect 47492 412632 47544 412684
rect 57888 412632 57940 412684
rect 204444 411884 204496 411936
rect 205732 411884 205784 411936
rect 358084 411884 358136 411936
rect 377036 411884 377088 411936
rect 48228 411272 48280 411324
rect 57888 411272 57940 411324
rect 217784 411272 217836 411324
rect 219256 411272 219308 411324
rect 3332 411204 3384 411256
rect 15844 411204 15896 411256
rect 205732 410524 205784 410576
rect 216772 410524 216824 410576
rect 216956 410524 217008 410576
rect 360016 410524 360068 410576
rect 377036 410524 377088 410576
rect 377496 410524 377548 410576
rect 50252 409844 50304 409896
rect 57888 409844 57940 409896
rect 377956 409844 378008 409896
rect 379428 409844 379480 409896
rect 359924 409096 359976 409148
rect 377404 409096 377456 409148
rect 50988 408484 51040 408536
rect 57888 408484 57940 408536
rect 576124 405628 576176 405680
rect 580172 405628 580224 405680
rect 199200 398216 199252 398268
rect 199752 398216 199804 398268
rect 198096 397808 198148 397860
rect 199108 397808 199160 397860
rect 520924 396720 520976 396772
rect 580356 396720 580408 396772
rect 44732 391892 44784 391944
rect 57060 391892 57112 391944
rect 209596 391892 209648 391944
rect 216680 391892 216732 391944
rect 359648 391892 359700 391944
rect 376944 391892 376996 391944
rect 207020 390464 207072 390516
rect 216680 390464 216732 390516
rect 358084 390464 358136 390516
rect 362960 390464 363012 390516
rect 376944 390464 376996 390516
rect 57520 389376 57572 389428
rect 52368 389104 52420 389156
rect 57244 389104 57296 389156
rect 57520 389104 57572 389156
rect 46112 389036 46164 389088
rect 57060 389036 57112 389088
rect 57520 388968 57572 389020
rect 206284 389172 206336 389224
rect 207020 389172 207072 389224
rect 200764 389104 200816 389156
rect 216680 389104 216732 389156
rect 359740 389104 359792 389156
rect 376944 389104 376996 389156
rect 57336 387744 57388 387796
rect 58624 387744 58676 387796
rect 58532 387676 58584 387728
rect 59360 387676 59412 387728
rect 57888 387132 57940 387184
rect 59728 387132 59780 387184
rect 56968 386316 57020 386368
rect 59728 386316 59780 386368
rect 369032 385704 369084 385756
rect 372804 385704 372856 385756
rect 219532 382372 219584 382424
rect 219900 382372 219952 382424
rect 217416 382236 217468 382288
rect 219532 382236 219584 382288
rect 57428 381624 57480 381676
rect 59544 381624 59596 381676
rect 197176 381488 197228 381540
rect 218244 381488 218296 381540
rect 55680 381012 55732 381064
rect 59452 381012 59504 381064
rect 196532 381012 196584 381064
rect 212816 381012 212868 381064
rect 196992 380944 197044 380996
rect 198188 380944 198240 380996
rect 199476 380944 199528 380996
rect 256056 380944 256108 380996
rect 55864 380876 55916 380928
rect 60096 380876 60148 380928
rect 143540 380876 143592 380928
rect 205916 380876 205968 380928
rect 375196 380876 375248 380928
rect 422852 380876 422904 380928
rect 47492 380808 47544 380860
rect 216864 380808 216916 380860
rect 48228 380740 48280 380792
rect 217324 380740 217376 380792
rect 52920 380672 52972 380724
rect 55864 380672 55916 380724
rect 50252 380604 50304 380656
rect 216956 380672 217008 380724
rect 367560 380672 367612 380724
rect 377956 380672 378008 380724
rect 160928 380604 160980 380656
rect 207388 380604 207440 380656
rect 365536 380604 365588 380656
rect 376668 380604 376720 380656
rect 377220 380604 377272 380656
rect 430948 380604 431000 380656
rect 146024 380536 146076 380588
rect 207296 380536 207348 380588
rect 360660 380536 360712 380588
rect 369860 380536 369912 380588
rect 371792 380536 371844 380588
rect 433616 380536 433668 380588
rect 59728 380468 59780 380520
rect 118424 380468 118476 380520
rect 133512 380468 133564 380520
rect 203156 380468 203208 380520
rect 204352 380468 204404 380520
rect 213644 380468 213696 380520
rect 358636 380468 358688 380520
rect 421104 380468 421156 380520
rect 57888 380400 57940 380452
rect 116032 380400 116084 380452
rect 135904 380400 135956 380452
rect 200580 380400 200632 380452
rect 202972 380400 203024 380452
rect 274640 380400 274692 380452
rect 369676 380400 369728 380452
rect 436008 380400 436060 380452
rect 48780 380332 48832 380384
rect 110972 380332 111024 380384
rect 131028 380332 131080 380384
rect 204628 380332 204680 380384
rect 262864 380332 262916 380384
rect 269764 380332 269816 380384
rect 366180 380332 366232 380384
rect 438492 380332 438544 380384
rect 58440 380264 58492 380316
rect 123484 380264 123536 380316
rect 163412 380264 163464 380316
rect 198004 380264 198056 380316
rect 200120 380264 200172 380316
rect 293960 380264 294012 380316
rect 363512 380264 363564 380316
rect 440884 380264 440936 380316
rect 58624 380196 58676 380248
rect 125968 380196 126020 380248
rect 128360 380196 128412 380248
rect 199292 380196 199344 380248
rect 200212 380196 200264 380248
rect 301504 380196 301556 380248
rect 360752 380196 360804 380248
rect 443460 380196 443512 380248
rect 45008 380128 45060 380180
rect 113548 380128 113600 380180
rect 121000 380128 121052 380180
rect 197912 380128 197964 380180
rect 201592 380128 201644 380180
rect 309048 380128 309100 380180
rect 362868 380128 362920 380180
rect 445944 380128 445996 380180
rect 155960 380060 156012 380112
rect 203248 380060 203300 380112
rect 158536 379992 158588 380044
rect 201868 379992 201920 380044
rect 214932 379992 214984 380044
rect 218060 379992 218112 380044
rect 165988 379924 166040 379976
rect 199016 379924 199068 379976
rect 213736 379924 213788 379976
rect 236000 379924 236052 379976
rect 240048 379924 240100 379976
rect 259460 379924 259512 379976
rect 207112 379856 207164 379908
rect 216496 379856 216548 379908
rect 243084 379856 243136 379908
rect 213644 379788 213696 379840
rect 237104 379788 237156 379840
rect 237380 379788 237432 379840
rect 265256 379788 265308 379840
rect 377404 379788 377456 379840
rect 377956 379788 378008 379840
rect 408684 379788 408736 379840
rect 212632 379720 212684 379772
rect 213920 379720 213972 379772
rect 220820 379720 220872 379772
rect 212724 379652 212776 379704
rect 219440 379652 219492 379704
rect 254492 379720 254544 379772
rect 369860 379720 369912 379772
rect 370964 379720 371016 379772
rect 413468 379720 413520 379772
rect 221004 379652 221056 379704
rect 255872 379652 255924 379704
rect 376484 379652 376536 379704
rect 376668 379652 376720 379704
rect 419448 379652 419500 379704
rect 208124 379584 208176 379636
rect 209504 379584 209556 379636
rect 216956 379584 217008 379636
rect 217784 379584 217836 379636
rect 218060 379584 218112 379636
rect 256976 379584 257028 379636
rect 375012 379584 375064 379636
rect 381176 379584 381228 379636
rect 426440 379584 426492 379636
rect 212540 379516 212592 379568
rect 258080 379516 258132 379568
rect 376576 379516 376628 379568
rect 434352 379516 434404 379568
rect 87696 379448 87748 379500
rect 209872 379448 209924 379500
rect 211344 379448 211396 379500
rect 213368 379448 213420 379500
rect 214104 379448 214156 379500
rect 219808 379448 219860 379500
rect 273260 379448 273312 379500
rect 274640 379448 274692 379500
rect 323308 379448 323360 379500
rect 325976 379448 326028 379500
rect 356612 379448 356664 379500
rect 364800 379448 364852 379500
rect 439044 379448 439096 379500
rect 59636 379380 59688 379432
rect 93492 379380 93544 379432
rect 202696 379380 202748 379432
rect 206928 379380 206980 379432
rect 268660 379380 268712 379432
rect 309048 379380 309100 379432
rect 315764 379380 315816 379432
rect 375380 379380 375432 379432
rect 435732 379380 435784 379432
rect 48872 379312 48924 379364
rect 88340 379312 88392 379364
rect 88800 379312 88852 379364
rect 209780 379312 209832 379364
rect 219624 379312 219676 379364
rect 219716 379312 219768 379364
rect 220268 379312 220320 379364
rect 271052 379312 271104 379364
rect 301504 379312 301556 379364
rect 313372 379312 313424 379364
rect 371148 379312 371200 379364
rect 375196 379312 375248 379364
rect 375288 379312 375340 379364
rect 408316 379312 408368 379364
rect 55956 379244 56008 379296
rect 90640 379244 90692 379296
rect 91376 379244 91428 379296
rect 211252 379244 211304 379296
rect 212540 379244 212592 379296
rect 212908 379244 212960 379296
rect 213368 379244 213420 379296
rect 253388 379244 253440 379296
rect 293960 379244 294012 379296
rect 310980 379244 311032 379296
rect 92388 379176 92440 379228
rect 201408 379176 201460 379228
rect 209872 379176 209924 379228
rect 219808 379176 219860 379228
rect 220728 379176 220780 379228
rect 46204 379108 46256 379160
rect 108212 379108 108264 379160
rect 114468 379108 114520 379160
rect 219900 379108 219952 379160
rect 220912 379108 220964 379160
rect 43996 379040 44048 379092
rect 105268 379040 105320 379092
rect 117136 379040 117188 379092
rect 44916 378972 44968 379024
rect 46204 378972 46256 379024
rect 50160 378972 50212 379024
rect 98460 378972 98512 379024
rect 112628 378972 112680 379024
rect 211252 379040 211304 379092
rect 221188 379040 221240 379092
rect 222016 379040 222068 379092
rect 57152 378904 57204 378956
rect 103520 378904 103572 378956
rect 55772 378836 55824 378888
rect 101036 378836 101088 378888
rect 44824 378768 44876 378820
rect 48872 378768 48924 378820
rect 90088 378768 90140 378820
rect 199016 378768 199068 378820
rect 209688 378972 209740 379024
rect 221004 378972 221056 379024
rect 208952 378904 209004 378956
rect 219716 378904 219768 378956
rect 201408 378836 201460 378888
rect 220820 378836 220872 378888
rect 222108 378836 222160 378888
rect 372436 378972 372488 379024
rect 380992 378972 381044 379024
rect 379796 378904 379848 378956
rect 397092 378904 397144 378956
rect 276940 378836 276992 378888
rect 361488 378836 361540 378888
rect 380900 378836 380952 378888
rect 205456 378768 205508 378820
rect 210332 378768 210384 378820
rect 212540 378768 212592 378820
rect 213460 378768 213512 378820
rect 219164 378768 219216 378820
rect 245384 378768 245436 378820
rect 359556 378768 359608 378820
rect 375472 378768 375524 378820
rect 379520 378768 379572 378820
rect 379980 378768 380032 378820
rect 403624 378768 403676 378820
rect 47860 378700 47912 378752
rect 96068 378700 96120 378752
rect 219716 378700 219768 378752
rect 219900 378700 219952 378752
rect 246028 378700 246080 378752
rect 375196 378700 375248 378752
rect 86592 378632 86644 378684
rect 208952 378632 209004 378684
rect 220728 378632 220780 378684
rect 247500 378632 247552 378684
rect 396080 378632 396132 378684
rect 199016 378564 199068 378616
rect 221280 378564 221332 378616
rect 250076 378564 250128 378616
rect 379336 378564 379388 378616
rect 379520 378564 379572 378616
rect 405832 378564 405884 378616
rect 219624 378496 219676 378548
rect 248604 378496 248656 378548
rect 380992 378496 381044 378548
rect 412364 378496 412416 378548
rect 108856 378428 108908 378480
rect 202696 378428 202748 378480
rect 210240 378428 210292 378480
rect 211344 378428 211396 378480
rect 222016 378428 222068 378480
rect 251180 378428 251232 378480
rect 380900 378428 380952 378480
rect 411260 378428 411312 378480
rect 113456 378360 113508 378412
rect 214104 378360 214156 378412
rect 222108 378360 222160 378412
rect 252284 378360 252336 378412
rect 343456 378360 343508 378412
rect 357532 378360 357584 378412
rect 358636 378360 358688 378412
rect 375472 378360 375524 378412
rect 376392 378360 376444 378412
rect 407580 378360 407632 378412
rect 111248 378292 111300 378344
rect 213368 378292 213420 378344
rect 220268 378292 220320 378344
rect 220912 378292 220964 378344
rect 274180 378292 274232 378344
rect 274272 378292 274324 378344
rect 302792 378292 302844 378344
rect 342260 378292 342312 378344
rect 343180 378292 343232 378344
rect 359372 378292 359424 378344
rect 48872 378224 48924 378276
rect 81440 378224 81492 378276
rect 93400 378224 93452 378276
rect 210240 378224 210292 378276
rect 210332 378224 210384 378276
rect 272064 378224 272116 378276
rect 277860 378224 277912 378276
rect 357440 378224 357492 378276
rect 377128 378292 377180 378344
rect 379428 378292 379480 378344
rect 426624 378292 426676 378344
rect 439044 378292 439096 378344
rect 516600 378292 516652 378344
rect 503076 378224 503128 378276
rect 517612 378224 517664 378276
rect 580264 378224 580316 378276
rect 46204 378156 46256 378208
rect 80428 378156 80480 378208
rect 85488 378156 85540 378208
rect 212540 378156 212592 378208
rect 274640 378156 274692 378208
rect 275652 378156 275704 378208
rect 356612 378156 356664 378208
rect 358636 378156 358688 378208
rect 503536 378156 503588 378208
rect 517704 378156 517756 378208
rect 580172 378156 580224 378208
rect 43260 378088 43312 378140
rect 199108 378088 199160 378140
rect 199844 378088 199896 378140
rect 201500 378088 201552 378140
rect 317420 378088 317472 378140
rect 357072 378088 357124 378140
rect 474832 378088 474884 378140
rect 54392 378020 54444 378072
rect 183192 378020 183244 378072
rect 198004 378020 198056 378072
rect 198832 378020 198884 378072
rect 300860 378020 300912 378072
rect 358728 378020 358780 378072
rect 460940 378020 460992 378072
rect 54300 377952 54352 378004
rect 182272 377952 182324 378004
rect 197452 377952 197504 378004
rect 298468 377952 298520 378004
rect 374368 377952 374420 378004
rect 458364 377952 458416 378004
rect 105544 377884 105596 377936
rect 215392 377884 215444 377936
rect 215760 377884 215812 377936
rect 217508 377884 217560 377936
rect 305828 377884 305880 377936
rect 370320 377884 370372 377936
rect 452752 377884 452804 377936
rect 150992 377816 151044 377868
rect 198096 377816 198148 377868
rect 198280 377816 198332 377868
rect 295892 377816 295944 377868
rect 365444 377816 365496 377868
rect 447508 377816 447560 377868
rect 148600 377748 148652 377800
rect 197268 377748 197320 377800
rect 197544 377748 197596 377800
rect 292672 377748 292724 377800
rect 373724 377748 373776 377800
rect 455604 377748 455656 377800
rect 196716 377680 196768 377732
rect 290924 377680 290976 377732
rect 196808 377612 196860 377664
rect 287704 377612 287756 377664
rect 359464 377612 359516 377664
rect 369860 377612 369912 377664
rect 196624 377544 196676 377596
rect 285956 377544 286008 377596
rect 368388 377544 368440 377596
rect 451004 377680 451056 377732
rect 98276 377476 98328 377528
rect 208952 377476 209004 377528
rect 212908 377476 212960 377528
rect 215760 377476 215812 377528
rect 219348 377476 219400 377528
rect 237380 377476 237432 377528
rect 369860 377476 369912 377528
rect 423404 377612 423456 377664
rect 372804 377544 372856 377596
rect 413100 377544 413152 377596
rect 379888 377476 379940 377528
rect 414572 377476 414624 377528
rect 199384 377408 199436 377460
rect 280712 377408 280764 377460
rect 367008 377408 367060 377460
rect 375288 377408 375340 377460
rect 197084 377340 197136 377392
rect 278044 377340 278096 377392
rect 415768 377408 415820 377460
rect 198740 377272 198792 377324
rect 274272 377272 274324 377324
rect 375288 377272 375340 377324
rect 377312 377272 377364 377324
rect 410064 377340 410116 377392
rect 153568 377204 153620 377256
rect 200396 377204 200448 377256
rect 373908 377204 373960 377256
rect 375932 377204 375984 377256
rect 402980 377272 403032 377324
rect 141056 377136 141108 377188
rect 200488 377136 200540 377188
rect 374460 377136 374512 377188
rect 379888 377136 379940 377188
rect 42156 377068 42208 377120
rect 199476 377068 199528 377120
rect 380900 376932 380952 376984
rect 381176 376932 381228 376984
rect 213000 376660 213052 376712
rect 283012 376660 283064 376712
rect 361304 376660 361356 376712
rect 477592 376660 477644 376712
rect 83464 376592 83516 376644
rect 207112 376592 207164 376644
rect 210148 376592 210200 376644
rect 320916 376592 320968 376644
rect 366272 376592 366324 376644
rect 480536 376592 480588 376644
rect 203892 376524 203944 376576
rect 273444 376524 273496 376576
rect 364156 376524 364208 376576
rect 473452 376524 473504 376576
rect 97172 376456 97224 376508
rect 211620 376456 211672 376508
rect 210056 376388 210108 376440
rect 212632 376388 212684 376440
rect 212540 376320 212592 376372
rect 213920 376456 213972 376508
rect 216404 376456 216456 376508
rect 217600 376456 217652 376508
rect 276020 376456 276072 376508
rect 362684 376456 362736 376508
rect 470876 376456 470928 376508
rect 213552 376388 213604 376440
rect 268108 376388 268160 376440
rect 364708 376388 364760 376440
rect 467932 376388 467984 376440
rect 138480 376252 138532 376304
rect 201776 376252 201828 376304
rect 213092 376320 213144 376372
rect 265900 376320 265952 376372
rect 367652 376320 367704 376372
rect 465080 376320 465132 376372
rect 263600 376252 263652 376304
rect 364248 376252 364300 376304
rect 427912 376252 427964 376304
rect 94688 376184 94740 376236
rect 212724 376184 212776 376236
rect 219256 376184 219308 376236
rect 270960 376184 271012 376236
rect 362776 376184 362828 376236
rect 425980 376184 426032 376236
rect 202512 376116 202564 376168
rect 248236 376116 248288 376168
rect 372528 376116 372580 376168
rect 418252 376116 418304 376168
rect 99472 376048 99524 376100
rect 213920 376048 213972 376100
rect 215852 376048 215904 376100
rect 260932 376048 260984 376100
rect 370412 376048 370464 376100
rect 416044 376048 416096 376100
rect 95976 375980 96028 376032
rect 213736 375980 213788 376032
rect 219532 375980 219584 376032
rect 258356 375980 258408 376032
rect 357164 375980 357216 376032
rect 208768 375912 208820 375964
rect 253572 375912 253624 375964
rect 379244 375980 379296 376032
rect 381176 375980 381228 376032
rect 436468 375980 436520 376032
rect 375840 375912 375892 375964
rect 416964 375912 417016 375964
rect 215024 375844 215076 375896
rect 250628 375844 250680 375896
rect 44640 375708 44692 375760
rect 216772 375776 216824 375828
rect 217600 375776 217652 375828
rect 104440 375640 104492 375692
rect 216588 375640 216640 375692
rect 217232 375640 217284 375692
rect 212540 375572 212592 375624
rect 214380 375572 214432 375624
rect 214932 375572 214984 375624
rect 216404 375572 216456 375624
rect 240048 375776 240100 375828
rect 213552 375368 213604 375420
rect 213736 375368 213788 375420
rect 107568 375300 107620 375352
rect 208308 375300 208360 375352
rect 217508 375300 217560 375352
rect 106464 375232 106516 375284
rect 208032 375232 208084 375284
rect 267556 375232 267608 375284
rect 102968 375164 103020 375216
rect 215300 375164 215352 375216
rect 216588 375164 216640 375216
rect 262772 375164 262824 375216
rect 101864 375096 101916 375148
rect 214472 375096 214524 375148
rect 261668 375096 261720 375148
rect 208124 375028 208176 375080
rect 279148 375028 279200 375080
rect 357164 375368 357216 375420
rect 368388 375368 368440 375420
rect 371240 375368 371292 375420
rect 372528 375368 372580 375420
rect 370228 375300 370280 375352
rect 431132 375300 431184 375352
rect 364064 375232 364116 375284
rect 377956 375232 378008 375284
rect 437756 375232 437808 375284
rect 369768 375164 369820 375216
rect 371792 375164 371844 375216
rect 373816 375164 373868 375216
rect 432236 375164 432288 375216
rect 372528 375096 372580 375148
rect 428280 375096 428332 375148
rect 364892 375028 364944 375080
rect 378140 375028 378192 375080
rect 379612 375028 379664 375080
rect 423956 375028 424008 375080
rect 85028 374960 85080 375012
rect 218152 374960 218204 375012
rect 218612 374960 218664 375012
rect 244280 374960 244332 375012
rect 368296 374960 368348 375012
rect 371516 374960 371568 375012
rect 372528 374960 372580 375012
rect 198004 374892 198056 374944
rect 342260 374892 342312 374944
rect 356888 374892 356940 374944
rect 372436 374892 372488 374944
rect 405372 374960 405424 375012
rect 361396 374824 361448 374876
rect 377220 374892 377272 374944
rect 418160 374892 418212 374944
rect 375656 374824 375708 374876
rect 378232 374824 378284 374876
rect 425152 374824 425204 374876
rect 357992 374756 358044 374808
rect 372988 374756 373040 374808
rect 421748 374756 421800 374808
rect 372528 374688 372580 374740
rect 419632 374688 419684 374740
rect 208032 374620 208084 374672
rect 219256 374620 219308 374672
rect 266360 374620 266412 374672
rect 377404 374620 377456 374672
rect 377956 374620 378008 374672
rect 371792 374552 371844 374604
rect 372528 374552 372580 374604
rect 429292 374620 429344 374672
rect 378140 374552 378192 374604
rect 379336 374552 379388 374604
rect 409972 374552 410024 374604
rect 359924 373260 359976 373312
rect 519360 373260 519412 373312
rect 519360 372580 519412 372632
rect 519636 372580 519688 372632
rect 359648 371832 359700 371884
rect 519176 371900 519228 371952
rect 519544 371900 519596 371952
rect 199476 370472 199528 370524
rect 359004 370472 359056 370524
rect 359004 369180 359056 369232
rect 359464 369180 359516 369232
rect 518992 369180 519044 369232
rect 199568 369112 199620 369164
rect 358912 369112 358964 369164
rect 359556 369112 359608 369164
rect 359556 366324 359608 366376
rect 519084 366324 519136 366376
rect 519360 366324 519412 366376
rect 199752 363604 199804 363656
rect 359096 363604 359148 363656
rect 519268 363604 519320 363656
rect 199568 362924 199620 362976
rect 199752 362924 199804 362976
rect 359188 362380 359240 362432
rect 359648 362380 359700 362432
rect 199752 362176 199804 362228
rect 359188 362176 359240 362228
rect 201408 360204 201460 360256
rect 206284 360204 206336 360256
rect 178684 360136 178736 360188
rect 196532 360136 196584 360188
rect 179880 360068 179932 360120
rect 197268 360068 197320 360120
rect 196532 359660 196584 359712
rect 197360 359660 197412 359712
rect 500776 359660 500828 359712
rect 517796 359592 517848 359644
rect 517980 359592 518032 359644
rect 339868 359524 339920 359576
rect 357072 359524 357124 359576
rect 498936 359524 498988 359576
rect 517888 359524 517940 359576
rect 190920 359456 190972 359508
rect 200764 359456 200816 359508
rect 201408 359456 201460 359508
rect 351736 359456 351788 359508
rect 358084 359456 358136 359508
rect 360200 359252 360252 359304
rect 361580 359252 361632 359304
rect 342260 358844 342312 358896
rect 357532 358844 357584 358896
rect 358636 358844 358688 358896
rect 338488 358776 338540 358828
rect 360200 358776 360252 358828
rect 510896 358776 510948 358828
rect 517520 358776 517572 358828
rect 218520 358708 218572 358760
rect 221188 358708 221240 358760
rect 378692 358708 378744 358760
rect 380900 358708 380952 358760
rect 215852 358640 215904 358692
rect 221004 358640 221056 358692
rect 219164 358504 219216 358556
rect 220820 358504 220872 358556
rect 217876 358232 217928 358284
rect 221280 358232 221332 358284
rect 379244 358232 379296 358284
rect 381084 358232 381136 358284
rect 214932 358164 214984 358216
rect 221096 358164 221148 358216
rect 54300 358028 54352 358080
rect 60096 358028 60148 358080
rect 182824 358028 182876 358080
rect 200120 358028 200172 358080
rect 342260 358028 342312 358080
rect 373816 358028 373868 358080
rect 381176 358028 381228 358080
rect 377036 357960 377088 358012
rect 380992 357960 381044 358012
rect 57152 357824 57204 357876
rect 59544 357824 59596 357876
rect 215760 357552 215812 357604
rect 220912 357552 220964 357604
rect 58532 356192 58584 356244
rect 59360 356192 59412 356244
rect 58624 355988 58676 356040
rect 59452 355988 59504 356040
rect 46296 303560 46348 303612
rect 57612 303560 57664 303612
rect 46388 300772 46440 300824
rect 57060 300772 57112 300824
rect 57428 300772 57480 300824
rect 57428 300636 57480 300688
rect 57612 300636 57664 300688
rect 520188 288396 520240 288448
rect 580264 288396 580316 288448
rect 519268 287036 519320 287088
rect 580356 287036 580408 287088
rect 200948 284248 201000 284300
rect 216680 284248 216732 284300
rect 361212 284248 361264 284300
rect 376944 284248 376996 284300
rect 203800 282820 203852 282872
rect 216864 282820 216916 282872
rect 366916 282820 366968 282872
rect 376760 282820 376812 282872
rect 55864 282684 55916 282736
rect 58440 282684 58492 282736
rect 52920 282344 52972 282396
rect 53196 282344 53248 282396
rect 54392 282140 54444 282192
rect 58716 282140 58768 282192
rect 200764 282140 200816 282192
rect 216680 282140 216732 282192
rect 358084 282140 358136 282192
rect 376944 282140 376996 282192
rect 58532 281460 58584 281512
rect 59728 281460 59780 281512
rect 212264 274728 212316 274780
rect 215668 274728 215720 274780
rect 213736 274660 213788 274712
rect 214104 274660 214156 274712
rect 215668 273912 215720 273964
rect 273168 273912 273220 273964
rect 43352 273572 43404 273624
rect 133420 273572 133472 273624
rect 45100 273504 45152 273556
rect 135904 273504 135956 273556
rect 219256 273504 219308 273556
rect 220820 273504 220872 273556
rect 266360 273504 266412 273556
rect 45468 273436 45520 273488
rect 138480 273436 138532 273488
rect 211712 273436 211764 273488
rect 214196 273436 214248 273488
rect 269764 273436 269816 273488
rect 370320 273436 370372 273488
rect 378140 273436 378192 273488
rect 378600 273436 378652 273488
rect 379520 273436 379572 273488
rect 427636 273436 427688 273488
rect 45192 273368 45244 273420
rect 140872 273368 140924 273420
rect 271144 273368 271196 273420
rect 374460 273368 374512 273420
rect 422852 273368 422904 273420
rect 45376 273300 45428 273352
rect 143540 273300 143592 273352
rect 213092 273300 213144 273352
rect 213368 273300 213420 273352
rect 213736 273300 213788 273352
rect 273260 273300 273312 273352
rect 366732 273300 366784 273352
rect 421104 273300 421156 273352
rect 45284 273232 45336 273284
rect 145932 273232 145984 273284
rect 206744 273232 206796 273284
rect 283472 273232 283524 273284
rect 370872 273232 370924 273284
rect 445944 273232 445996 273284
rect 42340 273164 42392 273216
rect 46020 273164 46072 273216
rect 378600 273164 378652 273216
rect 425244 273164 425296 273216
rect 212356 273096 212408 273148
rect 285956 273096 286008 273148
rect 369584 273096 369636 273148
rect 423404 273096 423456 273148
rect 209320 273028 209372 273080
rect 288164 273028 288216 273080
rect 356796 273028 356848 273080
rect 425980 273028 426032 273080
rect 216312 272960 216364 273012
rect 298468 272960 298520 273012
rect 358452 272960 358504 273012
rect 428188 272960 428240 273012
rect 210884 272892 210936 272944
rect 295892 272892 295944 272944
rect 372344 272892 372396 272944
rect 468484 272892 468536 272944
rect 42432 272824 42484 272876
rect 60832 272824 60884 272876
rect 202420 272824 202472 272876
rect 290924 272824 290976 272876
rect 373448 272824 373500 272876
rect 478420 272824 478472 272876
rect 48136 272756 48188 272808
rect 77116 272756 77168 272808
rect 203708 272756 203760 272808
rect 293316 272756 293368 272808
rect 363972 272756 364024 272808
rect 470876 272756 470928 272808
rect 50436 272688 50488 272740
rect 90732 272688 90784 272740
rect 207848 272688 207900 272740
rect 300860 272688 300912 272740
rect 365352 272688 365404 272740
rect 473452 272688 473504 272740
rect 48964 272620 49016 272672
rect 50252 272620 50304 272672
rect 51632 272620 51684 272672
rect 93676 272620 93728 272672
rect 205272 272620 205324 272672
rect 303436 272620 303488 272672
rect 368204 272620 368256 272672
rect 480812 272620 480864 272672
rect 48044 272552 48096 272604
rect 95884 272552 95936 272604
rect 206560 272552 206612 272604
rect 310980 272552 311032 272604
rect 362592 272552 362644 272604
rect 475844 272552 475896 272604
rect 50528 272484 50580 272536
rect 98460 272484 98512 272536
rect 107476 272484 107528 272536
rect 196900 272484 196952 272536
rect 200856 272484 200908 272536
rect 320916 272484 320968 272536
rect 361120 272484 361172 272536
rect 485964 272484 486016 272536
rect 49056 272416 49108 272468
rect 50068 272416 50120 272468
rect 46664 272348 46716 272400
rect 76012 272416 76064 272468
rect 58624 272348 58676 272400
rect 59452 272348 59504 272400
rect 62120 272348 62172 272400
rect 94412 272348 94464 272400
rect 50068 272280 50120 272332
rect 83004 272280 83056 272332
rect 374368 272280 374420 272332
rect 375104 272280 375156 272332
rect 58440 272212 58492 272264
rect 60740 272212 60792 272264
rect 100760 272212 100812 272264
rect 46480 272144 46532 272196
rect 51448 272144 51500 272196
rect 46572 272076 46624 272128
rect 48964 272076 49016 272128
rect 58716 272144 58768 272196
rect 60924 272144 60976 272196
rect 102140 272144 102192 272196
rect 95976 272076 96028 272128
rect 371792 272076 371844 272128
rect 373080 272076 373132 272128
rect 433340 272076 433392 272128
rect 52736 272008 52788 272060
rect 53288 272008 53340 272060
rect 60832 272008 60884 272060
rect 104900 272008 104952 272060
rect 373908 272008 373960 272060
rect 379612 272008 379664 272060
rect 396724 272008 396776 272060
rect 415860 272008 415912 272060
rect 48964 271940 49016 271992
rect 98000 271940 98052 271992
rect 370412 271940 370464 271992
rect 372344 271940 372396 271992
rect 430580 271940 430632 271992
rect 48228 271872 48280 271924
rect 107476 271872 107528 271924
rect 114468 271872 114520 271924
rect 127624 271872 127676 271924
rect 215852 271872 215904 271924
rect 216312 271872 216364 271924
rect 276020 271872 276072 271924
rect 356796 271872 356848 271924
rect 359372 271872 359424 271924
rect 43444 271804 43496 271856
rect 129740 271804 129792 271856
rect 154488 271804 154540 271856
rect 201684 271804 201736 271856
rect 343548 271804 343600 271856
rect 358636 271804 358688 271856
rect 360292 271872 360344 271924
rect 425704 271872 425756 271924
rect 427820 271872 427872 271924
rect 369492 271804 369544 271856
rect 458180 271804 458232 271856
rect 517704 271804 517756 271856
rect 517888 271804 517940 271856
rect 42248 271736 42300 271788
rect 123208 271736 123260 271788
rect 158628 271736 158680 271788
rect 205640 271736 205692 271788
rect 212172 271736 212224 271788
rect 307760 271736 307812 271788
rect 368020 271736 368072 271788
rect 455788 271736 455840 271788
rect 42524 271668 42576 271720
rect 52460 271668 52512 271720
rect 52828 271668 52880 271720
rect 54300 271668 54352 271720
rect 125600 271668 125652 271720
rect 151360 271668 151412 271720
rect 197636 271668 197688 271720
rect 202144 271668 202196 271720
rect 270500 271668 270552 271720
rect 363880 271668 363932 271720
rect 449900 271668 449952 271720
rect 57152 271600 57204 271652
rect 128360 271600 128412 271652
rect 157248 271600 157300 271652
rect 202880 271600 202932 271652
rect 214748 271600 214800 271652
rect 280160 271600 280212 271652
rect 370780 271600 370832 271652
rect 452660 271600 452712 271652
rect 54668 271532 54720 271584
rect 120080 271532 120132 271584
rect 161296 271532 161348 271584
rect 204260 271532 204312 271584
rect 216220 271532 216272 271584
rect 276020 271532 276072 271584
rect 368112 271532 368164 271584
rect 443000 271532 443052 271584
rect 53104 271464 53156 271516
rect 115940 271464 115992 271516
rect 164148 271464 164200 271516
rect 197728 271464 197780 271516
rect 205180 271464 205232 271516
rect 263600 271464 263652 271516
rect 372252 271464 372304 271516
rect 447140 271464 447192 271516
rect 46756 271396 46808 271448
rect 53840 271396 53892 271448
rect 54760 271396 54812 271448
rect 117320 271396 117372 271448
rect 166908 271396 166960 271448
rect 53196 271328 53248 271380
rect 113180 271328 113232 271380
rect 196624 271396 196676 271448
rect 197820 271396 197872 271448
rect 219072 271396 219124 271448
rect 277952 271396 278004 271448
rect 361028 271396 361080 271448
rect 426992 271396 427044 271448
rect 427084 271396 427136 271448
rect 432052 271396 432104 271448
rect 200304 271328 200356 271380
rect 203616 271328 203668 271380
rect 260840 271328 260892 271380
rect 362500 271328 362552 271380
rect 434720 271328 434772 271380
rect 503628 271328 503680 271380
rect 517612 271328 517664 271380
rect 51540 271260 51592 271312
rect 110420 271260 110472 271312
rect 197912 271260 197964 271312
rect 200120 271260 200172 271312
rect 210700 271260 210752 271312
rect 267832 271260 267884 271312
rect 343548 271260 343600 271312
rect 356796 271260 356848 271312
rect 366824 271260 366876 271312
rect 437480 271260 437532 271312
rect 52920 271192 52972 271244
rect 107660 271192 107712 271244
rect 183468 271192 183520 271244
rect 197452 271192 197504 271244
rect 198004 271192 198056 271244
rect 209412 271192 209464 271244
rect 264980 271192 265032 271244
rect 278688 271192 278740 271244
rect 357440 271192 357492 271244
rect 373632 271192 373684 271244
rect 440240 271192 440292 271244
rect 503628 271192 503680 271244
rect 517888 271192 517940 271244
rect 51816 271124 51868 271176
rect 104900 271124 104952 271176
rect 127624 271124 127676 271176
rect 196624 271124 196676 271176
rect 206652 271124 206704 271176
rect 258264 271124 258316 271176
rect 275928 271124 275980 271176
rect 356612 271124 356664 271176
rect 356796 271124 356848 271176
rect 358544 271124 358596 271176
rect 416044 271124 416096 271176
rect 426992 271124 427044 271176
rect 433340 271124 433392 271176
rect 440148 271124 440200 271176
rect 516600 271124 516652 271176
rect 51908 271056 51960 271108
rect 103520 271056 103572 271108
rect 209228 271056 209280 271108
rect 255320 271056 255372 271108
rect 379152 271056 379204 271108
rect 418160 271056 418212 271108
rect 50344 270988 50396 271040
rect 100760 270988 100812 271040
rect 210792 270988 210844 271040
rect 252560 270988 252612 271040
rect 374920 270988 374972 271040
rect 412732 270988 412784 271040
rect 54576 270920 54628 270972
rect 88340 270920 88392 270972
rect 214840 270920 214892 270972
rect 247040 270920 247092 270972
rect 374828 270920 374880 270972
rect 409880 270920 409932 270972
rect 213276 270852 213328 270904
rect 313280 270852 313332 270904
rect 183468 270512 183520 270564
rect 197728 270512 197780 270564
rect 197912 270512 197964 270564
rect 47952 270444 48004 270496
rect 147680 270444 147732 270496
rect 213000 270444 213052 270496
rect 213460 270444 213512 270496
rect 53196 270376 53248 270428
rect 86960 270376 87012 270428
rect 216864 270376 216916 270428
rect 219808 270444 219860 270496
rect 247040 270444 247092 270496
rect 280068 270444 280120 270496
rect 356612 270444 356664 270496
rect 357164 270444 357216 270496
rect 365536 270444 365588 270496
rect 368296 270444 368348 270496
rect 377220 270444 377272 270496
rect 377496 270444 377548 270496
rect 378508 270444 378560 270496
rect 379980 270444 380032 270496
rect 219900 270376 219952 270428
rect 220268 270376 220320 270428
rect 245660 270376 245712 270428
rect 378048 270376 378100 270428
rect 379244 270376 379296 270428
rect 411260 270444 411312 270496
rect 380440 270376 380492 270428
rect 407120 270376 407172 270428
rect 51724 270308 51776 270360
rect 84660 270308 84712 270360
rect 88248 270308 88300 270360
rect 109040 270308 109092 270360
rect 217876 270308 217928 270360
rect 249800 270308 249852 270360
rect 377956 270308 378008 270360
rect 408500 270308 408552 270360
rect 59728 270240 59780 270292
rect 61016 270240 61068 270292
rect 81440 270240 81492 270292
rect 111800 270240 111852 270292
rect 213460 270240 213512 270292
rect 244280 270240 244332 270292
rect 371608 270240 371660 270292
rect 373172 270240 373224 270292
rect 400220 270240 400272 270292
rect 52736 270172 52788 270224
rect 54576 270172 54628 270224
rect 85580 270172 85632 270224
rect 86868 270172 86920 270224
rect 110420 270172 110472 270224
rect 220636 270172 220688 270224
rect 248512 270172 248564 270224
rect 377036 270172 377088 270224
rect 378600 270172 378652 270224
rect 378692 270172 378744 270224
rect 401692 270172 401744 270224
rect 58624 270104 58676 270156
rect 89720 270104 89772 270156
rect 210332 270104 210384 270156
rect 213460 270104 213512 270156
rect 218428 270104 218480 270156
rect 218612 270104 218664 270156
rect 220728 270104 220780 270156
rect 251180 270104 251232 270156
rect 371056 270104 371108 270156
rect 59360 270036 59412 270088
rect 92480 270036 92532 270088
rect 210240 270036 210292 270088
rect 219716 270036 219768 270088
rect 252560 270036 252612 270088
rect 397460 270104 397512 270156
rect 379612 270036 379664 270088
rect 405740 270036 405792 270088
rect 54484 269968 54536 270020
rect 55956 269968 56008 270020
rect 88340 269968 88392 270020
rect 217232 269968 217284 270020
rect 218612 269968 218664 270020
rect 263600 269968 263652 270020
rect 374920 269968 374972 270020
rect 379796 269968 379848 270020
rect 379980 269968 380032 270020
rect 403624 269968 403676 270020
rect 80060 269900 80112 269952
rect 114560 269900 114612 269952
rect 219348 269900 219400 269952
rect 265164 269900 265216 269952
rect 368296 269900 368348 269952
rect 398840 269900 398892 269952
rect 57244 269832 57296 269884
rect 91100 269832 91152 269884
rect 113364 269832 113416 269884
rect 128360 269832 128412 269884
rect 219072 269832 219124 269884
rect 266360 269832 266412 269884
rect 378600 269832 378652 269884
rect 411352 269832 411404 269884
rect 61016 269764 61068 269816
rect 118700 269764 118752 269816
rect 213460 269764 213512 269816
rect 271880 269764 271932 269816
rect 370964 269764 371016 269816
rect 379980 269764 380032 269816
rect 413008 269764 413060 269816
rect 50620 269696 50672 269748
rect 54668 269696 54720 269748
rect 84200 269696 84252 269748
rect 208216 269696 208268 269748
rect 209412 269696 209464 269748
rect 237380 269696 237432 269748
rect 216588 269628 216640 269680
rect 262220 269628 262272 269680
rect 219164 269560 219216 269612
rect 219900 269560 219952 269612
rect 220728 269560 220780 269612
rect 218520 269492 218572 269544
rect 219256 269492 219308 269544
rect 251272 269560 251324 269612
rect 375748 269560 375800 269612
rect 376392 269560 376444 269612
rect 380440 269560 380492 269612
rect 218612 269356 218664 269408
rect 219072 269356 219124 269408
rect 218152 269288 218204 269340
rect 220268 269288 220320 269340
rect 214288 269220 214340 269272
rect 219624 269220 219676 269272
rect 220636 269220 220688 269272
rect 219348 269084 219400 269136
rect 219624 269084 219676 269136
rect 373632 269084 373684 269136
rect 375012 269152 375064 269204
rect 378692 269152 378744 269204
rect 377496 269084 377548 269136
rect 391940 269084 391992 269136
rect 47400 269016 47452 269068
rect 58624 269016 58676 269068
rect 128360 269016 128412 269068
rect 196992 269016 197044 269068
rect 208952 269016 209004 269068
rect 217232 269016 217284 269068
rect 258080 269016 258132 269068
rect 375840 269016 375892 269068
rect 416780 269016 416832 269068
rect 213644 268948 213696 269000
rect 215852 268948 215904 269000
rect 216220 268948 216272 269000
rect 216496 268948 216548 269000
rect 219440 268948 219492 269000
rect 253940 268948 253992 269000
rect 375656 268948 375708 269000
rect 375932 268948 375984 269000
rect 379888 268948 379940 269000
rect 414020 268948 414072 269000
rect 242900 268880 242952 268932
rect 388444 268880 388496 268932
rect 420920 268880 420972 268932
rect 214840 268812 214892 268864
rect 218428 268812 218480 268864
rect 244372 268812 244424 268864
rect 379152 268812 379204 268864
rect 409880 268812 409932 268864
rect 214380 268744 214432 268796
rect 218520 268744 218572 268796
rect 215852 268676 215904 268728
rect 236000 268744 236052 268796
rect 390560 268744 390612 268796
rect 419540 268744 419592 268796
rect 232504 268676 232556 268728
rect 259460 268676 259512 268728
rect 375932 268676 375984 268728
rect 402980 268676 403032 268728
rect 43628 268608 43680 268660
rect 46480 268608 46532 268660
rect 80060 268608 80112 268660
rect 213552 268608 213604 268660
rect 217048 268608 217100 268660
rect 217416 268608 217468 268660
rect 230480 268608 230532 268660
rect 259552 268608 259604 268660
rect 391940 268608 391992 268660
rect 418160 268608 418212 268660
rect 43812 268540 43864 268592
rect 46388 268540 46440 268592
rect 81440 268540 81492 268592
rect 229744 268540 229796 268592
rect 260840 268540 260892 268592
rect 43536 268472 43588 268524
rect 46204 268472 46256 268524
rect 86868 268472 86920 268524
rect 218520 268472 218572 268524
rect 256700 268472 256752 268524
rect 43720 268404 43772 268456
rect 46296 268404 46348 268456
rect 88248 268404 88300 268456
rect 217048 268404 217100 268456
rect 255320 268404 255372 268456
rect 47584 268336 47636 268388
rect 99380 268336 99432 268388
rect 202696 268336 202748 268388
rect 212172 268336 212224 268388
rect 268200 268336 268252 268388
rect 372436 268336 372488 268388
rect 374552 268336 374604 268388
rect 404360 268336 404412 268388
rect 43904 267656 43956 267708
rect 47584 267656 47636 267708
rect 371700 267656 371752 267708
rect 375196 267656 375248 267708
rect 434812 267656 434864 267708
rect 379060 267044 379112 267096
rect 437480 267044 437532 267096
rect 373816 266976 373868 267028
rect 375932 266976 375984 267028
rect 436100 266976 436152 267028
rect 219440 262896 219492 262948
rect 219716 262896 219768 262948
rect 340788 253852 340840 253904
rect 357072 253920 357124 253972
rect 357624 253920 357676 253972
rect 180156 253308 180208 253360
rect 197544 253308 197596 253360
rect 500868 253308 500920 253360
rect 517704 253308 517756 253360
rect 179328 253240 179380 253292
rect 197360 253240 197412 253292
rect 197636 253240 197688 253292
rect 339408 253240 339460 253292
rect 360200 253240 360252 253292
rect 499212 253240 499264 253292
rect 517796 253240 517848 253292
rect 191748 253172 191800 253224
rect 200764 253172 200816 253224
rect 351828 253172 351880 253224
rect 358084 253172 358136 253224
rect 517704 253172 517756 253224
rect 517980 253172 518032 253224
rect 510896 252560 510948 252612
rect 517520 252560 517572 252612
rect 58808 252492 58860 252544
rect 60924 252492 60976 252544
rect 214472 252492 214524 252544
rect 214748 252492 214800 252544
rect 218612 252492 218664 252544
rect 220820 252492 220872 252544
rect 56968 252424 57020 252476
rect 61016 252424 61068 252476
rect 215760 252424 215812 252476
rect 216404 252424 216456 252476
rect 232504 252492 232556 252544
rect 375288 252492 375340 252544
rect 377404 252492 377456 252544
rect 378416 252492 378468 252544
rect 434720 252492 434772 252544
rect 214748 252356 214800 252408
rect 229744 252424 229796 252476
rect 371792 252424 371844 252476
rect 373724 252424 373776 252476
rect 427084 252424 427136 252476
rect 375196 252356 375248 252408
rect 376576 252356 376628 252408
rect 377404 252356 377456 252408
rect 396724 252356 396776 252408
rect 378416 252288 378468 252340
rect 54484 251948 54536 252000
rect 60740 251948 60792 252000
rect 58532 251880 58584 251932
rect 106280 251880 106332 251932
rect 368388 251880 368440 251932
rect 372252 251880 372304 251932
rect 425704 251880 425756 251932
rect 53840 251812 53892 251864
rect 115940 251812 115992 251864
rect 216404 251812 216456 251864
rect 230480 251812 230532 251864
rect 375288 251812 375340 251864
rect 429200 251812 429252 251864
rect 58716 251608 58768 251660
rect 60832 251608 60884 251660
rect 46848 251132 46900 251184
rect 58532 251132 58584 251184
rect 372528 251132 372580 251184
rect 374828 251132 374880 251184
rect 375288 251132 375340 251184
rect 49148 251064 49200 251116
rect 53840 251064 53892 251116
rect 54300 251064 54352 251116
rect 519452 183540 519504 183592
rect 520188 183540 520240 183592
rect 580264 183540 580316 183592
rect 520096 183472 520148 183524
rect 580356 183472 580408 183524
rect 205088 177964 205140 178016
rect 216680 177964 216732 178016
rect 365260 177964 365312 178016
rect 376944 177964 376996 178016
rect 358084 175924 358136 175976
rect 376944 175924 376996 175976
rect 216680 175244 216732 175296
rect 200764 175176 200816 175228
rect 201500 175176 201552 175228
rect 207664 175176 207716 175228
rect 216956 175176 217008 175228
rect 363788 175176 363840 175228
rect 376944 175176 376996 175228
rect 50804 166948 50856 167000
rect 96068 166948 96120 167000
rect 374644 166948 374696 167000
rect 428280 166948 428332 167000
rect 49424 166880 49476 166932
rect 98460 166880 98512 166932
rect 376208 166880 376260 166932
rect 430948 166880 431000 166932
rect 50712 166812 50764 166864
rect 101036 166812 101088 166864
rect 358360 166812 358412 166864
rect 418436 166812 418488 166864
rect 53564 166744 53616 166796
rect 105820 166744 105872 166796
rect 212172 166744 212224 166796
rect 220820 166744 220872 166796
rect 358268 166744 358320 166796
rect 421012 166744 421064 166796
rect 52184 166676 52236 166728
rect 108212 166676 108264 166728
rect 210608 166676 210660 166728
rect 260932 166676 260984 166728
rect 356704 166676 356756 166728
rect 433616 166676 433668 166728
rect 59084 166608 59136 166660
rect 140872 166608 140924 166660
rect 204904 166608 204956 166660
rect 265900 166608 265952 166660
rect 372160 166608 372212 166660
rect 475844 166608 475896 166660
rect 56232 166540 56284 166592
rect 138480 166540 138532 166592
rect 204996 166540 205048 166592
rect 288256 166540 288308 166592
rect 370688 166540 370740 166592
rect 473452 166540 473504 166592
rect 59912 166472 59964 166524
rect 145932 166472 145984 166524
rect 206468 166472 206520 166524
rect 291016 166472 291068 166524
rect 373356 166472 373408 166524
rect 480904 166472 480956 166524
rect 59176 166404 59228 166456
rect 148508 166404 148560 166456
rect 202236 166404 202288 166456
rect 285956 166404 286008 166456
rect 365168 166404 365220 166456
rect 478420 166404 478472 166456
rect 58992 166336 59044 166388
rect 153292 166336 153344 166388
rect 209136 166336 209188 166388
rect 293316 166336 293368 166388
rect 367928 166336 367980 166388
rect 483388 166336 483440 166388
rect 41328 166268 41380 166320
rect 163320 166268 163372 166320
rect 211988 166268 212040 166320
rect 298468 166268 298520 166320
rect 366640 166268 366692 166320
rect 485964 166268 486016 166320
rect 54392 166200 54444 166252
rect 60740 166200 60792 166252
rect 369400 166200 369452 166252
rect 423404 166200 423456 166252
rect 357256 165792 357308 165844
rect 360292 165792 360344 165844
rect 46204 165656 46256 165708
rect 52184 165656 52236 165708
rect 111156 165656 111208 165708
rect 54300 165588 54352 165640
rect 116952 165588 117004 165640
rect 59820 165520 59872 165572
rect 150440 165520 150492 165572
rect 197360 165520 197412 165572
rect 197728 165520 197780 165572
rect 216036 165520 216088 165572
rect 325884 165520 325936 165572
rect 343272 165520 343324 165572
rect 356980 165588 357032 165640
rect 357532 165588 357584 165640
rect 375288 165588 375340 165640
rect 434352 165588 434404 165640
rect 362408 165520 362460 165572
rect 458364 165520 458416 165572
rect 56140 165452 56192 165504
rect 135260 165452 135312 165504
rect 210516 165452 210568 165504
rect 320916 165452 320968 165504
rect 360936 165452 360988 165504
rect 452660 165452 452712 165504
rect 55128 165384 55180 165436
rect 132500 165384 132552 165436
rect 213184 165384 213236 165436
rect 300860 165384 300912 165436
rect 369216 165384 369268 165436
rect 455420 165384 455472 165436
rect 54852 165316 54904 165368
rect 128360 165316 128412 165368
rect 214656 165316 214708 165368
rect 280160 165316 280212 165368
rect 363696 165316 363748 165368
rect 443460 165316 443512 165368
rect 56508 165248 56560 165300
rect 129740 165248 129792 165300
rect 211896 165248 211948 165300
rect 277400 165248 277452 165300
rect 370596 165248 370648 165300
rect 449900 165248 449952 165300
rect 56324 165180 56376 165232
rect 125876 165180 125928 165232
rect 218980 165180 219032 165232
rect 283380 165180 283432 165232
rect 372068 165180 372120 165232
rect 447324 165180 447376 165232
rect 55036 165112 55088 165164
rect 123484 165112 123536 165164
rect 183468 165112 183520 165164
rect 197360 165112 197412 165164
rect 206376 165112 206428 165164
rect 267740 165112 267792 165164
rect 373264 165112 373316 165164
rect 445852 165112 445904 165164
rect 503260 165112 503312 165164
rect 517612 165112 517664 165164
rect 56048 165044 56100 165096
rect 120908 165044 120960 165096
rect 218888 165044 218940 165096
rect 276020 165044 276072 165096
rect 366548 165044 366600 165096
rect 438492 165044 438544 165096
rect 440148 165044 440200 165096
rect 516600 165044 516652 165096
rect 52092 164976 52144 165028
rect 115940 164976 115992 165028
rect 183192 164976 183244 165028
rect 197452 164976 197504 165028
rect 216128 164976 216180 165028
rect 273444 164976 273496 165028
rect 367836 164976 367888 165028
rect 435916 164976 435968 165028
rect 503352 164976 503404 165028
rect 517888 164976 517940 165028
rect 54944 164908 54996 164960
rect 113548 164908 113600 164960
rect 114652 164908 114704 164960
rect 196716 164908 196768 164960
rect 202328 164908 202380 164960
rect 255320 164908 255372 164960
rect 374736 164908 374788 164960
rect 440884 164908 440936 164960
rect 510528 164908 510580 164960
rect 517520 164908 517572 164960
rect 52000 164840 52052 164892
rect 91744 164840 91796 164892
rect 114468 164840 114520 164892
rect 114744 164840 114796 164892
rect 196624 164840 196676 164892
rect 203524 164840 203576 164892
rect 249800 164840 249852 164892
rect 343456 164840 343508 164892
rect 356704 164840 356756 164892
rect 357256 164840 357308 164892
rect 365076 164840 365128 164892
rect 412640 164840 412692 164892
rect 53472 164772 53524 164824
rect 94596 164772 94648 164824
rect 94780 164772 94832 164824
rect 118148 164772 118200 164824
rect 215944 164772 215996 164824
rect 258080 164772 258132 164824
rect 378876 164772 378928 164824
rect 416044 164772 416096 164824
rect 50896 164704 50948 164756
rect 89996 164704 90048 164756
rect 211804 164704 211856 164756
rect 252560 164704 252612 164756
rect 376116 164704 376168 164756
rect 409880 164704 409932 164756
rect 56416 164636 56468 164688
rect 88340 164636 88392 164688
rect 91744 164636 91796 164688
rect 103520 164636 103572 164688
rect 214564 164636 214616 164688
rect 247040 164636 247092 164688
rect 378968 164636 379020 164688
rect 407120 164636 407172 164688
rect 98644 164296 98696 164348
rect 100760 164296 100812 164348
rect 427820 164296 427872 164348
rect 435088 164296 435140 164348
rect 100024 164228 100076 164280
rect 103520 164228 103572 164280
rect 58532 164160 58584 164212
rect 59912 164160 59964 164212
rect 57520 164092 57572 164144
rect 117872 164160 117924 164212
rect 219624 164160 219676 164212
rect 264980 164160 265032 164212
rect 374828 164160 374880 164212
rect 429660 164160 429712 164212
rect 56968 163956 57020 164008
rect 59452 163956 59504 164008
rect 53656 163888 53708 163940
rect 110972 164092 111024 164144
rect 218336 164092 218388 164144
rect 219072 164092 219124 164144
rect 263784 164092 263836 164144
rect 374460 164092 374512 164144
rect 376116 164092 376168 164144
rect 379704 164092 379756 164144
rect 426440 164092 426492 164144
rect 213368 164024 213420 164076
rect 236092 164024 236144 164076
rect 379520 164024 379572 164076
rect 426532 164024 426584 164076
rect 374920 163956 374972 164008
rect 396172 163956 396224 164008
rect 212264 163888 212316 163940
rect 213368 163888 213420 163940
rect 374368 163888 374420 163940
rect 396080 163888 396132 163940
rect 51448 163820 51500 163872
rect 57060 163820 57112 163872
rect 95240 163820 95292 163872
rect 50160 163752 50212 163804
rect 56508 163752 56560 163804
rect 96620 163752 96672 163804
rect 48964 163684 49016 163736
rect 55036 163684 55088 163736
rect 98000 163684 98052 163736
rect 59912 163616 59964 163668
rect 106372 163616 106424 163668
rect 46296 163548 46348 163600
rect 53656 163548 53708 163600
rect 109316 163548 109368 163600
rect 376116 163548 376168 163600
rect 422300 163548 422352 163600
rect 59452 163480 59504 163532
rect 118884 163480 118936 163532
rect 213368 163480 213420 163532
rect 273812 163480 273864 163532
rect 371792 163480 371844 163532
rect 374920 163480 374972 163532
rect 432236 163480 432288 163532
rect 46480 162800 46532 162852
rect 50896 162800 50948 162852
rect 217048 162800 217100 162852
rect 217876 162800 217928 162852
rect 218520 162800 218572 162852
rect 218980 162800 219032 162852
rect 46388 162732 46440 162784
rect 52092 162732 52144 162784
rect 214748 162732 214800 162784
rect 260840 162800 260892 162852
rect 371700 162800 371752 162852
rect 372528 162800 372580 162852
rect 375932 162800 375984 162852
rect 376576 162800 376628 162852
rect 377496 162800 377548 162852
rect 379612 162800 379664 162852
rect 379796 162800 379848 162852
rect 436192 162800 436244 162852
rect 219348 162732 219400 162784
rect 259460 162732 259512 162784
rect 375840 162732 375892 162784
rect 378968 162732 379020 162784
rect 379060 162732 379112 162784
rect 437940 162732 437992 162784
rect 216404 162664 216456 162716
rect 259552 162664 259604 162716
rect 372528 162664 372580 162716
rect 427820 162664 427872 162716
rect 217324 162596 217376 162648
rect 258172 162596 258224 162648
rect 376300 162596 376352 162648
rect 418712 162596 418764 162648
rect 376484 162528 376536 162580
rect 379244 162528 379296 162580
rect 419540 162528 419592 162580
rect 376576 162460 376628 162512
rect 379796 162460 379848 162512
rect 214656 162392 214708 162444
rect 215760 162392 215812 162444
rect 219348 162392 219400 162444
rect 379612 162256 379664 162308
rect 418160 162256 418212 162308
rect 52092 162188 52144 162240
rect 112076 162188 112128 162240
rect 373540 162188 373592 162240
rect 376208 162188 376260 162240
rect 420920 162188 420972 162240
rect 50896 162120 50948 162172
rect 115756 162120 115808 162172
rect 219164 161780 219216 161832
rect 266360 162120 266412 162172
rect 372344 162120 372396 162172
rect 375012 162120 375064 162172
rect 430580 162120 430632 162172
rect 219532 161780 219584 161832
rect 218980 161508 219032 161560
rect 236644 161508 236696 161560
rect 217876 161440 217928 161492
rect 235264 161440 235316 161492
rect 378968 161440 379020 161492
rect 396724 161440 396776 161492
rect 58716 148996 58768 149048
rect 106280 148996 106332 149048
rect 213552 148996 213604 149048
rect 274732 148996 274784 149048
rect 373816 148996 373868 149048
rect 401600 148996 401652 149048
rect 216312 148928 216364 148980
rect 277400 148928 277452 148980
rect 371608 148928 371660 148980
rect 372436 148928 372488 148980
rect 400220 148928 400272 148980
rect 46572 148792 46624 148844
rect 54944 148792 54996 148844
rect 80060 148792 80112 148844
rect 47860 148724 47912 148776
rect 53472 148724 53524 148776
rect 78680 148724 78732 148776
rect 49056 148656 49108 148708
rect 52000 148656 52052 148708
rect 81440 148656 81492 148708
rect 52920 148588 52972 148640
rect 55864 148588 55916 148640
rect 100024 148588 100076 148640
rect 213276 148588 213328 148640
rect 238760 148588 238812 148640
rect 46112 148520 46164 148572
rect 59820 148520 59872 148572
rect 107660 148520 107712 148572
rect 214932 148520 214984 148572
rect 240140 148520 240192 148572
rect 59176 148452 59228 148504
rect 107752 148452 107804 148504
rect 213736 148452 213788 148504
rect 241520 148452 241572 148504
rect 374736 148452 374788 148504
rect 397460 148452 397512 148504
rect 53564 148384 53616 148436
rect 114652 148384 114704 148436
rect 213092 148384 213144 148436
rect 215024 148384 215076 148436
rect 270500 148384 270552 148436
rect 374828 148384 374880 148436
rect 398840 148384 398892 148436
rect 53104 148316 53156 148368
rect 114744 148316 114796 148368
rect 213460 148316 213512 148368
rect 215944 148316 215996 148368
rect 271880 148316 271932 148368
rect 373080 148316 373132 148368
rect 375196 148316 375248 148368
rect 434720 148316 434772 148368
rect 48228 147568 48280 147620
rect 58900 147568 58952 147620
rect 59176 147568 59228 147620
rect 210884 147568 210936 147620
rect 214564 147568 214616 147620
rect 214932 147568 214984 147620
rect 371056 147568 371108 147620
rect 374736 147568 374788 147620
rect 212356 147500 212408 147552
rect 213276 147500 213328 147552
rect 368296 147500 368348 147552
rect 374828 147500 374880 147552
rect 208308 147432 208360 147484
rect 213184 147432 213236 147484
rect 213736 147432 213788 147484
rect 48044 146208 48096 146260
rect 51724 146208 51776 146260
rect 56968 146208 57020 146260
rect 57244 146208 57296 146260
rect 59084 146208 59136 146260
rect 59360 146208 59412 146260
rect 213736 146276 213788 146328
rect 91100 146208 91152 146260
rect 179052 146208 179104 146260
rect 197636 146208 197688 146260
rect 53196 146140 53248 146192
rect 86960 146140 87012 146192
rect 179696 146140 179748 146192
rect 197544 146140 197596 146192
rect 214472 146140 214524 146192
rect 215852 146140 215904 146192
rect 236000 146208 236052 146260
rect 236644 146208 236696 146260
rect 256700 146208 256752 146260
rect 274824 146208 274876 146260
rect 356796 146208 356848 146260
rect 377588 146208 377640 146260
rect 378048 146208 378100 146260
rect 378600 146208 378652 146260
rect 379336 146208 379388 146260
rect 235264 146140 235316 146192
rect 255412 146140 255464 146192
rect 338488 146140 338540 146192
rect 360200 146140 360252 146192
rect 377404 146140 377456 146192
rect 377956 146140 378008 146192
rect 403072 146208 403124 146260
rect 58624 146072 58676 146124
rect 59176 146072 59228 146124
rect 59728 146072 59780 146124
rect 60740 146072 60792 146124
rect 66260 146072 66312 146124
rect 59360 146004 59412 146056
rect 92480 146072 92532 146124
rect 219256 146072 219308 146124
rect 251180 146072 251232 146124
rect 340236 146072 340288 146124
rect 357624 146072 357676 146124
rect 375932 146072 375984 146124
rect 378508 146072 378560 146124
rect 396724 146140 396776 146192
rect 416780 146140 416832 146192
rect 500224 146140 500276 146192
rect 517520 146140 517572 146192
rect 517704 146140 517756 146192
rect 379244 146072 379296 146124
rect 379980 146072 380032 146124
rect 412640 146072 412692 146124
rect 498660 146072 498712 146124
rect 517796 146072 517848 146124
rect 66444 146004 66496 146056
rect 93860 146004 93912 146056
rect 215760 146004 215812 146056
rect 217968 146004 218020 146056
rect 249892 146004 249944 146056
rect 379336 146004 379388 146056
rect 411260 146004 411312 146056
rect 56140 145936 56192 145988
rect 88432 145936 88484 145988
rect 218428 145936 218480 145988
rect 219808 145936 219860 145988
rect 219900 145936 219952 145988
rect 59176 145868 59228 145920
rect 89812 145868 89864 145920
rect 217048 145868 217100 145920
rect 251272 145936 251324 145988
rect 377956 145936 378008 145988
rect 378048 145936 378100 145988
rect 379152 145936 379204 145988
rect 409972 145936 410024 145988
rect 224224 145868 224276 145920
rect 244280 145868 244332 145920
rect 374552 145868 374604 145920
rect 374828 145868 374880 145920
rect 408500 145868 408552 145920
rect 54576 145800 54628 145852
rect 54852 145800 54904 145852
rect 85580 145800 85632 145852
rect 216128 145800 216180 145852
rect 216864 145800 216916 145852
rect 247132 145800 247184 145852
rect 404360 145800 404412 145852
rect 58716 145732 58768 145784
rect 84200 145732 84252 145784
rect 218152 145732 218204 145784
rect 218888 145732 218940 145784
rect 245660 145732 245712 145784
rect 374552 145732 374604 145784
rect 375656 145732 375708 145784
rect 402980 145732 403032 145784
rect 56416 145664 56468 145716
rect 84292 145664 84344 145716
rect 216220 145664 216272 145716
rect 216496 145664 216548 145716
rect 242900 145664 242952 145716
rect 378784 145664 378836 145716
rect 407212 145664 407264 145716
rect 50068 145596 50120 145648
rect 54392 145596 54444 145648
rect 82820 145596 82872 145648
rect 214840 145596 214892 145648
rect 224224 145596 224276 145648
rect 224316 145596 224368 145648
rect 244372 145596 244424 145648
rect 376392 145596 376444 145648
rect 405740 145596 405792 145648
rect 517520 145596 517572 145648
rect 580264 145596 580316 145648
rect 58624 145528 58676 145580
rect 91192 145528 91244 145580
rect 191288 145528 191340 145580
rect 201500 145528 201552 145580
rect 204904 145528 204956 145580
rect 216956 145528 217008 145580
rect 248420 145528 248472 145580
rect 280068 145528 280120 145580
rect 307668 145528 307720 145580
rect 351644 145528 351696 145580
rect 358084 145528 358136 145580
rect 358728 145528 358780 145580
rect 510528 145528 510580 145580
rect 517796 145528 517848 145580
rect 580356 145528 580408 145580
rect 51724 145460 51776 145512
rect 77300 145460 77352 145512
rect 218520 145460 218572 145512
rect 236092 145460 236144 145512
rect 378692 145460 378744 145512
rect 396080 145460 396132 145512
rect 48136 145392 48188 145444
rect 54484 145392 54536 145444
rect 75920 145392 75972 145444
rect 219716 145392 219768 145444
rect 253940 145392 253992 145444
rect 378876 145392 378928 145444
rect 396172 145392 396224 145444
rect 46664 145324 46716 145376
rect 54760 145324 54812 145376
rect 76012 145324 76064 145376
rect 219808 145324 219860 145376
rect 252652 145324 252704 145376
rect 379888 145324 379940 145376
rect 414020 145324 414072 145376
rect 377588 145256 377640 145308
rect 411352 145256 411404 145308
rect 216036 144984 216088 145036
rect 224316 144984 224368 145036
rect 54668 144848 54720 144900
rect 56048 144848 56100 144900
rect 56416 144848 56468 144900
rect 214288 144848 214340 144900
rect 216956 144848 217008 144900
rect 217140 144848 217192 144900
rect 307668 144848 307720 144900
rect 356612 144848 356664 144900
rect 51816 144780 51868 144832
rect 58716 144780 58768 144832
rect 209412 144780 209464 144832
rect 213460 144780 213512 144832
rect 373908 144780 373960 144832
rect 376024 144780 376076 144832
rect 376392 144780 376444 144832
rect 53288 144712 53340 144764
rect 58624 144712 58676 144764
rect 213000 144712 213052 144764
rect 216036 144712 216088 144764
rect 377404 144916 377456 144968
rect 47584 144644 47636 144696
rect 55956 144644 56008 144696
rect 56324 144644 56376 144696
rect 376392 144644 376444 144696
rect 56232 144576 56284 144628
rect 375748 144576 375800 144628
rect 378784 144576 378836 144628
rect 56324 144372 56376 144424
rect 3516 97928 3568 97980
rect 21364 97928 21416 97980
rect 520188 79976 520240 80028
rect 580448 79976 580500 80028
rect 42616 70320 42668 70372
rect 57612 70320 57664 70372
rect 209044 70320 209096 70372
rect 216680 70320 216732 70372
rect 362316 70320 362368 70372
rect 376944 70320 376996 70372
rect 358728 68280 358780 68332
rect 376944 68280 376996 68332
rect 358084 68144 358136 68196
rect 358728 68144 358780 68196
rect 204904 67600 204956 67652
rect 216680 67600 216732 67652
rect 54484 59712 54536 59764
rect 77116 59712 77168 59764
rect 378876 59712 378928 59764
rect 397092 59712 397144 59764
rect 54392 59644 54444 59696
rect 83096 59644 83148 59696
rect 218520 59644 218572 59696
rect 236000 59644 236052 59696
rect 378692 59644 378744 59696
rect 396080 59644 396132 59696
rect 58992 59576 59044 59628
rect 100760 59576 100812 59628
rect 214472 59576 214524 59628
rect 237104 59576 237156 59628
rect 374552 59576 374604 59628
rect 403072 59576 403124 59628
rect 54576 59508 54628 59560
rect 101772 59508 101824 59560
rect 217876 59508 217928 59560
rect 255872 59508 255924 59560
rect 378968 59508 379020 59560
rect 416964 59508 417016 59560
rect 58900 59440 58952 59492
rect 107568 59440 107620 59492
rect 218980 59440 219032 59492
rect 256976 59440 257028 59492
rect 377496 59440 377548 59492
rect 423956 59440 424008 59492
rect 52276 59372 52328 59424
rect 113548 59372 113600 59424
rect 216588 59372 216640 59424
rect 262864 59372 262916 59424
rect 376116 59372 376168 59424
rect 422852 59372 422904 59424
rect 56048 59304 56100 59356
rect 84200 59304 84252 59356
rect 217968 59304 218020 59356
rect 358084 59304 358136 59356
rect 379888 59304 379940 59356
rect 414572 59304 414624 59356
rect 59728 59236 59780 59288
rect 94504 59236 94556 59288
rect 379612 59236 379664 59288
rect 418160 59236 418212 59288
rect 57060 59168 57112 59220
rect 95884 59168 95936 59220
rect 214656 59168 214708 59220
rect 259460 59168 259512 59220
rect 371884 59168 371936 59220
rect 410708 59168 410760 59220
rect 56508 59100 56560 59152
rect 96988 59100 97040 59152
rect 214748 59100 214800 59152
rect 261668 59100 261720 59152
rect 279240 59100 279292 59152
rect 356612 59100 356664 59152
rect 376300 59100 376352 59152
rect 419356 59100 419408 59152
rect 55036 59032 55088 59084
rect 98092 59032 98144 59084
rect 205548 59032 205600 59084
rect 290924 59032 290976 59084
rect 376484 59032 376536 59084
rect 420644 59032 420696 59084
rect 56324 58964 56376 59016
rect 102784 58964 102836 59016
rect 213828 58964 213880 59016
rect 300860 58964 300912 59016
rect 376208 58964 376260 59016
rect 421748 58964 421800 59016
rect 55864 58896 55916 58948
rect 103888 58896 103940 58948
rect 212448 58896 212500 58948
rect 315856 58896 315908 58948
rect 360844 58896 360896 58948
rect 416044 58896 416096 58948
rect 59820 58828 59872 58880
rect 108672 58828 108724 58880
rect 202788 58828 202840 58880
rect 308496 58828 308548 58880
rect 358176 58828 358228 58880
rect 423496 58828 423548 58880
rect 49608 58760 49660 58812
rect 110972 58760 111024 58812
rect 209596 58760 209648 58812
rect 320916 58760 320968 58812
rect 366456 58760 366508 58812
rect 468484 58760 468536 58812
rect 50988 58692 51040 58744
rect 148508 58692 148560 58744
rect 209504 58692 209556 58744
rect 325884 58692 325936 58744
rect 363604 58692 363656 58744
rect 475844 58692 475896 58744
rect 53012 58624 53064 58676
rect 150900 58624 150952 58676
rect 219072 58624 219124 58676
rect 428188 58624 428240 58676
rect 216404 58556 216456 58608
rect 260656 58556 260708 58608
rect 375932 58556 375984 58608
rect 404176 58556 404228 58608
rect 57888 57876 57940 57928
rect 204904 57876 204956 57928
rect 211068 57876 211120 57928
rect 323308 57876 323360 57928
rect 343180 57876 343232 57928
rect 357532 57876 357584 57928
rect 376668 57876 376720 57928
rect 485964 57876 486016 57928
rect 503260 57876 503312 57928
rect 517612 57876 517664 57928
rect 51632 57808 51684 57860
rect 145564 57808 145616 57860
rect 183284 57808 183336 57860
rect 197452 57808 197504 57860
rect 206192 57808 206244 57860
rect 313372 57808 313424 57860
rect 343456 57808 343508 57860
rect 356704 57808 356756 57860
rect 365628 57808 365680 57860
rect 470876 57808 470928 57860
rect 503536 57808 503588 57860
rect 517888 57808 517940 57860
rect 43996 57740 44048 57792
rect 123484 57740 123536 57792
rect 183468 57740 183520 57792
rect 197360 57740 197412 57792
rect 218244 57740 218296 57792
rect 318248 57740 318300 57792
rect 379428 57740 379480 57792
rect 478420 57740 478472 57792
rect 53748 57672 53800 57724
rect 133420 57672 133472 57724
rect 215116 57672 215168 57724
rect 310980 57672 311032 57724
rect 367744 57672 367796 57724
rect 465908 57672 465960 57724
rect 52368 57604 52420 57656
rect 130844 57604 130896 57656
rect 208676 57604 208728 57656
rect 303436 57604 303488 57656
rect 371148 57604 371200 57656
rect 460940 57604 460992 57656
rect 54208 57536 54260 57588
rect 128360 57536 128412 57588
rect 215668 57536 215720 57588
rect 305828 57536 305880 57588
rect 369124 57536 369176 57588
rect 445852 57536 445904 57588
rect 44088 57468 44140 57520
rect 57244 57468 57296 57520
rect 57888 57468 57940 57520
rect 115940 57468 115992 57520
rect 210976 57468 211028 57520
rect 295892 57468 295944 57520
rect 362224 57468 362276 57520
rect 438492 57468 438544 57520
rect 60004 57400 60056 57452
rect 125876 57400 125928 57452
rect 210424 57400 210476 57452
rect 293316 57400 293368 57452
rect 364984 57400 365036 57452
rect 433524 57400 433576 57452
rect 55956 57332 56008 57384
rect 99380 57332 99432 57384
rect 218796 57332 218848 57384
rect 298100 57332 298152 57384
rect 371976 57332 372028 57384
rect 435916 57332 435968 57384
rect 59268 57264 59320 57316
rect 93584 57264 93636 57316
rect 215208 57264 215260 57316
rect 287612 57264 287664 57316
rect 370504 57264 370556 57316
rect 430948 57264 431000 57316
rect 51724 57196 51776 57248
rect 78220 57196 78272 57248
rect 218704 57196 218756 57248
rect 258356 57196 258408 57248
rect 378416 57196 378468 57248
rect 415492 57196 415544 57248
rect 54760 57128 54812 57180
rect 76012 57128 76064 57180
rect 54300 56516 54352 56568
rect 116676 56516 116728 56568
rect 219992 56516 220044 56568
rect 408316 56516 408368 56568
rect 53104 56448 53156 56500
rect 113824 56448 113876 56500
rect 213552 56448 213604 56500
rect 273260 56448 273312 56500
rect 376576 56448 376628 56500
rect 436376 56448 436428 56500
rect 52092 56380 52144 56432
rect 112076 56380 112128 56432
rect 216312 56380 216364 56432
rect 276940 56380 276992 56432
rect 375288 56380 375340 56432
rect 434628 56380 434680 56432
rect 53656 56312 53708 56364
rect 109500 56312 109552 56364
rect 215024 56312 215076 56364
rect 271052 56312 271104 56364
rect 374920 56312 374972 56364
rect 432236 56312 432288 56364
rect 42708 56244 42760 56296
rect 90732 56244 90784 56296
rect 219900 56244 219952 56296
rect 268476 56244 268528 56296
rect 379244 56244 379296 56296
rect 412640 56244 412692 56296
rect 58624 56176 58676 56228
rect 92204 56176 92256 56228
rect 218612 56176 218664 56228
rect 266360 56176 266412 56228
rect 376392 56176 376444 56228
rect 408684 56176 408736 56228
rect 56416 56108 56468 56160
rect 88708 56108 88760 56160
rect 215760 56108 215812 56160
rect 250076 56108 250128 56160
rect 379336 56108 379388 56160
rect 411260 56108 411312 56160
rect 54852 56040 54904 56092
rect 86500 56040 86552 56092
rect 217048 56040 217100 56092
rect 251916 56040 251968 56092
rect 373816 56040 373868 56092
rect 401692 56040 401744 56092
rect 52000 55972 52052 56024
rect 81900 55972 81952 56024
rect 216128 55972 216180 56024
rect 247684 55972 247736 56024
rect 374736 55972 374788 56024
rect 399484 55972 399536 56024
rect 58716 55904 58768 55956
rect 85396 55904 85448 55956
rect 216036 55904 216088 55956
rect 245292 55904 245344 55956
rect 53472 55836 53524 55888
rect 79508 55836 79560 55888
rect 213276 55836 213328 55888
rect 239220 55836 239272 55888
rect 213184 55768 213236 55820
rect 241612 55768 241664 55820
rect 50896 55156 50948 55208
rect 114560 55156 114612 55208
rect 218888 55156 218940 55208
rect 245660 55156 245712 55208
rect 378784 55156 378836 55208
rect 407212 55156 407264 55208
rect 53564 55088 53616 55140
rect 113272 55088 113324 55140
rect 215944 55088 215996 55140
rect 271880 55088 271932 55140
rect 379060 55088 379112 55140
rect 437480 55088 437532 55140
rect 52184 55020 52236 55072
rect 110420 55020 110472 55072
rect 219532 55020 219584 55072
rect 266452 55020 266504 55072
rect 375196 55020 375248 55072
rect 433432 55020 433484 55072
rect 59912 54952 59964 55004
rect 106280 54952 106332 55004
rect 219624 54952 219676 55004
rect 264980 54952 265032 55004
rect 375012 54952 375064 55004
rect 430580 54952 430632 55004
rect 56968 54884 57020 54936
rect 91192 54884 91244 54936
rect 218336 54884 218388 54936
rect 263600 54884 263652 54936
rect 375104 54884 375156 54936
rect 429200 54884 429252 54936
rect 53196 54816 53248 54868
rect 86960 54816 87012 54868
rect 219716 54816 219768 54868
rect 253940 54816 253992 54868
rect 379796 54816 379848 54868
rect 426440 54816 426492 54868
rect 59084 54748 59136 54800
rect 92480 54748 92532 54800
rect 218428 54748 218480 54800
rect 252560 54748 252612 54800
rect 379520 54748 379572 54800
rect 426532 54748 426584 54800
rect 59176 54680 59228 54732
rect 89812 54680 89864 54732
rect 219256 54680 219308 54732
rect 251180 54680 251232 54732
rect 377588 54680 377640 54732
rect 411352 54680 411404 54732
rect 54944 54612 54996 54664
rect 80060 54612 80112 54664
rect 217140 54612 217192 54664
rect 248420 54612 248472 54664
rect 378048 54612 378100 54664
rect 409880 54612 409932 54664
rect 214840 54544 214892 54596
rect 244372 54544 244424 54596
rect 376024 54544 376076 54596
rect 405832 54544 405884 54596
rect 216496 54476 216548 54528
rect 242900 54476 242952 54528
rect 374828 54476 374880 54528
rect 404360 54476 404412 54528
rect 213368 54408 213420 54460
rect 273352 54408 273404 54460
rect 372528 54408 372580 54460
rect 434720 54408 434772 54460
rect 213460 54340 213512 54392
rect 237380 54340 237432 54392
rect 374644 54340 374696 54392
rect 397460 54340 397512 54392
rect 214564 54272 214616 54324
rect 240140 54272 240192 54324
rect 372436 54272 372488 54324
rect 400220 54272 400272 54324
rect 3424 20612 3476 20664
rect 10324 20612 10376 20664
rect 572 3408 624 3460
rect 57244 3408 57296 3460
rect 125876 3408 125928 3460
rect 366364 3408 366416 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 638246 3464 684247
rect 3424 638240 3476 638246
rect 3424 638182 3476 638188
rect 40052 636886 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 57796 700324 57848 700330
rect 57796 700266 57848 700272
rect 40040 636880 40092 636886
rect 40040 636822 40092 636828
rect 56508 633684 56560 633690
rect 56508 633626 56560 633632
rect 55036 633616 55088 633622
rect 55036 633558 55088 633564
rect 54852 633480 54904 633486
rect 54852 633422 54904 633428
rect 3516 632868 3568 632874
rect 3516 632810 3568 632816
rect 3424 632460 3476 632466
rect 3424 632402 3476 632408
rect 3436 632097 3464 632402
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 568546 3464 579935
rect 3424 568540 3476 568546
rect 3424 568482 3476 568488
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3422 482216 3478 482225
rect 3422 482151 3478 482160
rect 3332 411256 3384 411262
rect 3332 411198 3384 411204
rect 3344 410553 3372 411198
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3436 58585 3464 482151
rect 3528 306241 3556 632810
rect 3608 632800 3660 632806
rect 3608 632742 3660 632748
rect 3620 358465 3648 632742
rect 54864 568002 54892 633422
rect 54944 630760 54996 630766
rect 54944 630702 54996 630708
rect 54852 567996 54904 568002
rect 54852 567938 54904 567944
rect 10324 563712 10376 563718
rect 10324 563654 10376 563660
rect 3700 480956 3752 480962
rect 3700 480898 3752 480904
rect 3712 462641 3740 480898
rect 3698 462632 3754 462641
rect 3698 462567 3754 462576
rect 3606 358456 3662 358465
rect 3606 358391 3662 358400
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 10336 20670 10364 563654
rect 21364 554804 21416 554810
rect 21364 554746 21416 554752
rect 11704 514820 11756 514826
rect 11704 514762 11756 514768
rect 11716 488102 11744 514762
rect 11704 488096 11756 488102
rect 11704 488038 11756 488044
rect 15844 486464 15896 486470
rect 15844 486406 15896 486412
rect 15856 411262 15884 486406
rect 15844 411256 15896 411262
rect 15844 411198 15896 411204
rect 21376 97986 21404 554746
rect 54956 550458 54984 630702
rect 54944 550452 54996 550458
rect 54944 550394 54996 550400
rect 55048 550254 55076 633558
rect 55128 633548 55180 633554
rect 55128 633490 55180 633496
rect 55140 550526 55168 633490
rect 56416 631032 56468 631038
rect 56416 630974 56468 630980
rect 56324 630964 56376 630970
rect 56324 630906 56376 630912
rect 55128 550520 55180 550526
rect 55128 550462 55180 550468
rect 55036 550248 55088 550254
rect 55036 550190 55088 550196
rect 56336 550050 56364 630906
rect 56428 550186 56456 630974
rect 56520 550322 56548 633626
rect 57704 630828 57756 630834
rect 57704 630770 57756 630776
rect 57610 628688 57666 628697
rect 57610 628623 57666 628632
rect 57426 622432 57482 622441
rect 57426 622367 57482 622376
rect 57334 597952 57390 597961
rect 57334 597887 57390 597896
rect 57242 591832 57298 591841
rect 57242 591767 57298 591776
rect 57150 589112 57206 589121
rect 57150 589047 57206 589056
rect 57058 582992 57114 583001
rect 57058 582927 57114 582936
rect 57072 566778 57100 582927
rect 57164 569226 57192 589047
rect 57152 569220 57204 569226
rect 57152 569162 57204 569168
rect 57060 566772 57112 566778
rect 57060 566714 57112 566720
rect 57256 559706 57284 591767
rect 57348 568478 57376 597887
rect 57440 591394 57468 622367
rect 57518 619712 57574 619721
rect 57518 619647 57574 619656
rect 57428 591388 57480 591394
rect 57428 591330 57480 591336
rect 57426 579728 57482 579737
rect 57426 579663 57482 579672
rect 57336 568472 57388 568478
rect 57336 568414 57388 568420
rect 57244 559700 57296 559706
rect 57244 559642 57296 559648
rect 57440 556986 57468 579663
rect 57532 566642 57560 619647
rect 57520 566636 57572 566642
rect 57520 566578 57572 566584
rect 57428 556980 57480 556986
rect 57428 556922 57480 556928
rect 57624 551342 57652 628623
rect 57612 551336 57664 551342
rect 57612 551278 57664 551284
rect 56508 550316 56560 550322
rect 56508 550258 56560 550264
rect 56416 550180 56468 550186
rect 56416 550122 56468 550128
rect 57716 550118 57744 630770
rect 57808 607617 57836 700266
rect 104912 639606 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 170324 700398 170352 703520
rect 235184 700466 235212 703520
rect 235172 700460 235224 700466
rect 235172 700402 235224 700408
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 147588 683188 147640 683194
rect 147588 683130 147640 683136
rect 104900 639600 104952 639606
rect 104900 639542 104952 639548
rect 144920 634160 144972 634166
rect 144920 634102 144972 634108
rect 109960 634024 110012 634030
rect 109960 633966 110012 633972
rect 120908 634024 120960 634030
rect 120908 633966 120960 633972
rect 86776 633888 86828 633894
rect 86776 633830 86828 633836
rect 77300 633684 77352 633690
rect 77300 633626 77352 633632
rect 65524 631032 65576 631038
rect 77312 630986 77340 633626
rect 80244 633616 80296 633622
rect 80244 633558 80296 633564
rect 80256 630986 80284 633558
rect 86788 630986 86816 633830
rect 106648 633752 106700 633758
rect 106648 633694 106700 633700
rect 104072 633684 104124 633690
rect 104072 633626 104124 633632
rect 100668 633616 100720 633622
rect 100668 633558 100720 633564
rect 91836 633548 91888 633554
rect 91836 633490 91888 633496
rect 95056 633548 95108 633554
rect 95056 633490 95108 633496
rect 88708 633480 88760 633486
rect 88708 633422 88760 633428
rect 65576 630980 65826 630986
rect 65524 630974 65826 630980
rect 65536 630958 65826 630974
rect 71240 630970 71622 630986
rect 71228 630964 71622 630970
rect 71280 630958 71622 630964
rect 77312 630958 77418 630986
rect 80256 630958 80638 630986
rect 83214 630970 83504 630986
rect 83214 630964 83516 630970
rect 83214 630958 83464 630964
rect 71228 630906 71280 630912
rect 86434 630958 86816 630986
rect 88720 630986 88748 633422
rect 91848 630986 91876 633490
rect 95068 630986 95096 633490
rect 100680 630986 100708 633558
rect 104084 630986 104112 633626
rect 106660 630986 106688 633694
rect 109972 630986 110000 633966
rect 112536 633956 112588 633962
rect 112536 633898 112588 633904
rect 112548 630986 112576 633898
rect 115664 633820 115716 633826
rect 115664 633762 115716 633768
rect 115676 630986 115704 633762
rect 88720 630958 89010 630986
rect 91848 630958 92230 630986
rect 94806 630958 95096 630986
rect 100602 630958 100708 630986
rect 103822 630958 104112 630986
rect 106398 630958 106688 630986
rect 109618 630958 110000 630986
rect 112194 630958 112576 630986
rect 115414 630958 115704 630986
rect 83464 630906 83516 630912
rect 59360 630896 59412 630902
rect 97908 630896 97960 630902
rect 59360 630838 59412 630844
rect 57888 630692 57940 630698
rect 57888 630634 57940 630640
rect 57794 607608 57850 607617
rect 57794 607543 57850 607552
rect 57900 604081 57928 630634
rect 59266 625832 59322 625841
rect 59266 625767 59322 625776
rect 58990 616312 59046 616321
rect 58990 616247 59046 616256
rect 57886 604072 57942 604081
rect 57886 604007 57942 604016
rect 57794 595232 57850 595241
rect 57794 595167 57850 595176
rect 57808 581670 57836 595167
rect 57796 581664 57848 581670
rect 57796 581606 57848 581612
rect 57794 573472 57850 573481
rect 57794 573407 57850 573416
rect 57808 554198 57836 573407
rect 57796 554192 57848 554198
rect 57796 554134 57848 554140
rect 57704 550112 57756 550118
rect 57704 550054 57756 550060
rect 56324 550044 56376 550050
rect 56324 549986 56376 549992
rect 57900 517993 57928 604007
rect 58898 601352 58954 601361
rect 58898 601287 58954 601296
rect 58624 591388 58676 591394
rect 58624 591330 58676 591336
rect 58530 576872 58586 576881
rect 58530 576807 58586 576816
rect 58544 566574 58572 576807
rect 58532 566568 58584 566574
rect 58532 566510 58584 566516
rect 58636 549914 58664 591330
rect 58806 585712 58862 585721
rect 58806 585647 58862 585656
rect 58716 581664 58768 581670
rect 58716 581606 58768 581612
rect 58728 550390 58756 581606
rect 58820 568138 58848 585647
rect 58808 568132 58860 568138
rect 58808 568074 58860 568080
rect 58912 563854 58940 601287
rect 59004 568070 59032 616247
rect 59174 613592 59230 613601
rect 59174 613527 59230 613536
rect 59082 610192 59138 610201
rect 59082 610127 59138 610136
rect 58992 568064 59044 568070
rect 58992 568006 59044 568012
rect 58900 563848 58952 563854
rect 58900 563790 58952 563796
rect 59096 556850 59124 610127
rect 59084 556844 59136 556850
rect 59084 556786 59136 556792
rect 59188 555490 59216 613527
rect 59280 561134 59308 625767
rect 59268 561128 59320 561134
rect 59268 561070 59320 561076
rect 59176 555484 59228 555490
rect 59176 555426 59228 555432
rect 59372 552786 59400 630838
rect 74644 630834 74842 630850
rect 97960 630844 98026 630850
rect 97908 630838 98026 630844
rect 74632 630828 74842 630834
rect 74684 630822 74842 630828
rect 97920 630822 98026 630838
rect 74632 630770 74684 630776
rect 62948 630760 63000 630766
rect 69296 630760 69348 630766
rect 63000 630708 63250 630714
rect 62948 630702 63250 630708
rect 62960 630686 63250 630702
rect 69046 630708 69296 630714
rect 69046 630702 69348 630708
rect 69046 630686 69336 630702
rect 59464 630414 60030 630442
rect 117990 630426 118188 630442
rect 117990 630420 118200 630426
rect 117990 630414 118148 630420
rect 59464 562426 59492 630414
rect 120566 630414 120764 630442
rect 118148 630362 118200 630368
rect 59542 570788 59598 570797
rect 59542 570723 59598 570732
rect 59452 562420 59504 562426
rect 59452 562362 59504 562368
rect 59556 558210 59584 570723
rect 59912 569220 59964 569226
rect 59912 569162 59964 569168
rect 59544 558204 59596 558210
rect 59544 558146 59596 558152
rect 59924 557534 59952 569162
rect 60740 568472 60792 568478
rect 60740 568414 60792 568420
rect 113180 568472 113232 568478
rect 113180 568414 113232 568420
rect 60030 568126 60320 568154
rect 60292 565214 60320 568126
rect 60280 565208 60332 565214
rect 60280 565150 60332 565156
rect 60752 557534 60780 568414
rect 106280 568404 106332 568410
rect 106280 568346 106332 568352
rect 99564 568336 99616 568342
rect 99564 568278 99616 568284
rect 96712 568268 96764 568274
rect 96712 568210 96764 568216
rect 87052 568200 87104 568206
rect 62606 568126 62896 568154
rect 62120 566772 62172 566778
rect 62120 566714 62172 566720
rect 62132 557534 62160 566714
rect 62868 565146 62896 568126
rect 64984 568126 65182 568154
rect 67640 568132 67692 568138
rect 63500 567860 63552 567866
rect 63500 567802 63552 567808
rect 62856 565140 62908 565146
rect 62856 565082 62908 565088
rect 59924 557506 60412 557534
rect 60752 557506 60964 557534
rect 62132 557506 62436 557534
rect 59372 552758 60320 552786
rect 58716 550384 58768 550390
rect 58716 550326 58768 550332
rect 58624 549908 58676 549914
rect 58624 549850 58676 549856
rect 60292 547963 60320 552758
rect 60384 549982 60412 557506
rect 60372 549976 60424 549982
rect 60372 549918 60424 549924
rect 60936 547963 60964 557506
rect 61660 549364 61712 549370
rect 61660 549306 61712 549312
rect 61672 547963 61700 549306
rect 62408 547963 62436 557506
rect 63132 554124 63184 554130
rect 63132 554066 63184 554072
rect 63144 547963 63172 554066
rect 63512 552786 63540 567802
rect 64880 566500 64932 566506
rect 64880 566442 64932 566448
rect 63592 560992 63644 560998
rect 63592 560934 63644 560940
rect 63604 557534 63632 560934
rect 63604 557506 64552 557534
rect 63512 552758 63816 552786
rect 63788 547963 63816 552758
rect 64524 547963 64552 557506
rect 64892 549250 64920 566442
rect 64984 549370 65012 568126
rect 68402 568126 68784 568154
rect 70978 568126 71360 568154
rect 67640 568074 67692 568080
rect 66352 567928 66404 567934
rect 66352 567870 66404 567876
rect 65064 559564 65116 559570
rect 65064 559506 65116 559512
rect 65076 557534 65104 559506
rect 66364 557534 66392 567870
rect 65076 557506 66024 557534
rect 66364 557506 66760 557534
rect 64972 549364 65024 549370
rect 64972 549306 65024 549312
rect 64892 549222 65288 549250
rect 65260 547963 65288 549222
rect 65996 547963 66024 557506
rect 66732 547963 66760 557506
rect 67652 552770 67680 568074
rect 68756 562494 68784 568126
rect 71332 565282 71360 568126
rect 73816 568126 74198 568154
rect 76774 568126 77064 568154
rect 71320 565276 71372 565282
rect 71320 565218 71372 565224
rect 73816 564466 73844 568126
rect 74540 568064 74592 568070
rect 74540 568006 74592 568012
rect 71780 564460 71832 564466
rect 71780 564402 71832 564408
rect 73804 564460 73856 564466
rect 73804 564402 73856 564408
rect 69020 563780 69072 563786
rect 69020 563722 69072 563728
rect 68744 562488 68796 562494
rect 68744 562430 68796 562436
rect 69032 552770 69060 563722
rect 69112 562352 69164 562358
rect 69112 562294 69164 562300
rect 69124 557534 69152 562294
rect 70400 561060 70452 561066
rect 70400 561002 70452 561008
rect 70412 557534 70440 561002
rect 71792 557534 71820 564402
rect 69124 557506 69612 557534
rect 70412 557506 70992 557534
rect 71792 557506 72464 557534
rect 67640 552764 67692 552770
rect 67640 552706 67692 552712
rect 68836 552764 68888 552770
rect 68836 552706 68888 552712
rect 69020 552764 69072 552770
rect 69020 552706 69072 552712
rect 68098 552664 68154 552673
rect 68098 552599 68154 552608
rect 67364 550520 67416 550526
rect 67364 550462 67416 550468
rect 67376 547963 67404 550462
rect 68112 547963 68140 552599
rect 68848 547963 68876 552706
rect 69584 547963 69612 557506
rect 70308 552764 70360 552770
rect 70308 552706 70360 552712
rect 70320 547963 70348 552706
rect 70964 547963 70992 557506
rect 71688 554056 71740 554062
rect 71688 553998 71740 554004
rect 71700 547963 71728 553998
rect 72436 547963 72464 557506
rect 73160 555620 73212 555626
rect 73160 555562 73212 555568
rect 73172 547963 73200 555562
rect 73804 550044 73856 550050
rect 73804 549986 73856 549992
rect 73816 547963 73844 549986
rect 74552 547963 74580 568006
rect 74632 565480 74684 565486
rect 74632 565422 74684 565428
rect 74644 557534 74672 565422
rect 77036 565418 77064 568126
rect 79888 568126 79994 568154
rect 82570 568126 82768 568154
rect 85790 568126 86080 568154
rect 87052 568142 87104 568148
rect 78680 567996 78732 568002
rect 78680 567938 78732 567944
rect 77024 565412 77076 565418
rect 77024 565354 77076 565360
rect 75920 562420 75972 562426
rect 75920 562362 75972 562368
rect 75932 557534 75960 562362
rect 74644 557506 75316 557534
rect 75932 557506 76052 557534
rect 75288 547963 75316 557506
rect 76024 547963 76052 557506
rect 78692 552770 78720 567938
rect 79888 565350 79916 568126
rect 82740 565554 82768 568126
rect 82912 566636 82964 566642
rect 82912 566578 82964 566584
rect 84200 566636 84252 566642
rect 84200 566578 84252 566584
rect 82728 565548 82780 565554
rect 82728 565490 82780 565496
rect 79876 565344 79928 565350
rect 79876 565286 79928 565292
rect 78772 562420 78824 562426
rect 78772 562362 78824 562368
rect 78784 557534 78812 562362
rect 80060 558272 80112 558278
rect 80060 558214 80112 558220
rect 80072 557534 80100 558214
rect 82924 557534 82952 566578
rect 84212 557534 84240 566578
rect 86052 565418 86080 568126
rect 86960 567996 87012 568002
rect 86960 567938 87012 567944
rect 84844 565412 84896 565418
rect 84844 565354 84896 565360
rect 86040 565412 86092 565418
rect 86040 565354 86092 565360
rect 78784 557506 78904 557534
rect 80072 557506 80376 557534
rect 82924 557506 83228 557534
rect 84212 557506 84608 557534
rect 78680 552764 78732 552770
rect 78680 552706 78732 552712
rect 76748 552696 76800 552702
rect 76748 552638 76800 552644
rect 76760 547963 76788 552638
rect 77392 551336 77444 551342
rect 77392 551278 77444 551284
rect 77404 547963 77432 551278
rect 78128 550044 78180 550050
rect 78128 549986 78180 549992
rect 78140 547963 78168 549986
rect 78876 547963 78904 557506
rect 79600 552764 79652 552770
rect 79600 552706 79652 552712
rect 79612 547963 79640 552706
rect 80348 547963 80376 557506
rect 80980 557048 81032 557054
rect 80980 556990 81032 556996
rect 80992 547963 81020 556990
rect 81716 556980 81768 556986
rect 81716 556922 81768 556928
rect 81728 547963 81756 556922
rect 82452 552764 82504 552770
rect 82452 552706 82504 552712
rect 82464 547963 82492 552706
rect 83200 547963 83228 557506
rect 83924 550316 83976 550322
rect 83924 550258 83976 550264
rect 83936 547963 83964 550258
rect 84580 547963 84608 557506
rect 84856 550594 84884 565354
rect 85672 559632 85724 559638
rect 85672 559574 85724 559580
rect 85684 557534 85712 559574
rect 85684 557506 86080 557534
rect 84844 550588 84896 550594
rect 84844 550530 84896 550536
rect 85304 550316 85356 550322
rect 85304 550258 85356 550264
rect 85316 547963 85344 550258
rect 86052 547963 86080 557506
rect 86972 552786 87000 567938
rect 87064 557534 87092 568142
rect 88366 568126 88472 568154
rect 88444 559774 88472 568126
rect 91112 568126 91586 568154
rect 93860 568132 93912 568138
rect 89720 565548 89772 565554
rect 89720 565490 89772 565496
rect 88432 559768 88484 559774
rect 88432 559710 88484 559716
rect 88432 558408 88484 558414
rect 88432 558350 88484 558356
rect 87064 557506 88196 557534
rect 86972 552758 87460 552786
rect 86776 550588 86828 550594
rect 86776 550530 86828 550536
rect 86788 547963 86816 550530
rect 87432 547963 87460 552758
rect 88168 547963 88196 557506
rect 88444 552838 88472 558350
rect 88432 552832 88484 552838
rect 88432 552774 88484 552780
rect 89628 552832 89680 552838
rect 89628 552774 89680 552780
rect 89732 552786 89760 565490
rect 89812 559700 89864 559706
rect 89812 559642 89864 559648
rect 89824 552906 89852 559642
rect 89812 552900 89864 552906
rect 89812 552842 89864 552848
rect 91008 552900 91060 552906
rect 91008 552842 91060 552848
rect 88892 550452 88944 550458
rect 88892 550394 88944 550400
rect 88904 547963 88932 550394
rect 89640 547963 89668 552774
rect 89732 552758 90404 552786
rect 90376 547963 90404 552758
rect 91020 547963 91048 552842
rect 91112 550458 91140 568126
rect 94162 568126 94544 568154
rect 93860 568074 93912 568080
rect 91192 563848 91244 563854
rect 91192 563790 91244 563796
rect 91204 557534 91232 563790
rect 92572 561128 92624 561134
rect 92572 561070 92624 561076
rect 91204 557506 91784 557534
rect 91100 550452 91152 550458
rect 91100 550394 91152 550400
rect 91756 547963 91784 557506
rect 92584 548162 92612 561070
rect 93872 557534 93900 568074
rect 94516 564942 94544 568126
rect 94504 564936 94556 564942
rect 94504 564878 94556 564884
rect 96724 557534 96752 568210
rect 97000 568126 97382 568154
rect 97000 565486 97028 568126
rect 98092 568064 98144 568070
rect 98092 568006 98144 568012
rect 96988 565480 97040 565486
rect 96988 565422 97040 565428
rect 98104 557534 98132 568006
rect 98644 558340 98696 558346
rect 98644 558282 98696 558288
rect 93872 557506 93992 557534
rect 96724 557506 97488 557534
rect 98104 557506 98224 557534
rect 93216 550248 93268 550254
rect 93216 550190 93268 550196
rect 92508 548134 92612 548162
rect 92508 547944 92536 548134
rect 93228 547963 93256 550190
rect 93964 547963 93992 557506
rect 94596 551336 94648 551342
rect 94596 551278 94648 551284
rect 94608 547963 94636 551278
rect 96068 550588 96120 550594
rect 96068 550530 96120 550536
rect 95332 550384 95384 550390
rect 95332 550326 95384 550332
rect 95344 547963 95372 550326
rect 96080 547963 96108 550530
rect 96804 550452 96856 550458
rect 96804 550394 96856 550400
rect 96816 547963 96844 550394
rect 97460 547963 97488 557506
rect 98196 547963 98224 557506
rect 98656 550594 98684 558282
rect 99576 557534 99604 568278
rect 99958 568126 100248 568154
rect 100220 565486 100248 568126
rect 102888 568126 103178 568154
rect 104912 568126 105754 568154
rect 100208 565480 100260 565486
rect 100208 565422 100260 565428
rect 102784 564936 102836 564942
rect 102784 564878 102836 564884
rect 100760 564460 100812 564466
rect 100760 564402 100812 564408
rect 99576 557506 100432 557534
rect 98644 550588 98696 550594
rect 98644 550530 98696 550536
rect 98920 550180 98972 550186
rect 98920 550122 98972 550128
rect 98932 547963 98960 550122
rect 99656 550112 99708 550118
rect 99656 550054 99708 550060
rect 99668 547963 99696 550054
rect 100404 547963 100432 557506
rect 100772 552838 100800 564402
rect 100852 558204 100904 558210
rect 100852 558146 100904 558152
rect 100864 557534 100892 558146
rect 100864 557506 101076 557534
rect 100760 552832 100812 552838
rect 100760 552774 100812 552780
rect 101048 547963 101076 557506
rect 102508 556844 102560 556850
rect 102508 556786 102560 556792
rect 101772 552832 101824 552838
rect 101772 552774 101824 552780
rect 101784 547963 101812 552774
rect 102520 547963 102548 556786
rect 102796 550186 102824 564878
rect 102888 564466 102916 568126
rect 104164 565208 104216 565214
rect 104164 565150 104216 565156
rect 102876 564460 102928 564466
rect 102876 564402 102928 564408
rect 103520 559768 103572 559774
rect 103520 559710 103572 559716
rect 103244 554192 103296 554198
rect 103244 554134 103296 554140
rect 102784 550180 102836 550186
rect 102784 550122 102836 550128
rect 103256 547963 103284 554134
rect 103532 550474 103560 559710
rect 104176 550594 104204 565150
rect 104912 558414 104940 568126
rect 104900 558408 104952 558414
rect 104900 558350 104952 558356
rect 106292 552702 106320 568346
rect 107672 568126 108974 568154
rect 110616 568126 111550 568154
rect 106924 562488 106976 562494
rect 106924 562430 106976 562436
rect 106280 552696 106332 552702
rect 106280 552638 106332 552644
rect 104164 550588 104216 550594
rect 104164 550530 104216 550536
rect 105360 550588 105412 550594
rect 105360 550530 105412 550536
rect 103532 550446 104664 550474
rect 103980 550112 104032 550118
rect 103980 550054 104032 550060
rect 103992 547963 104020 550054
rect 104636 547963 104664 550446
rect 105372 547963 105400 550530
rect 106936 550526 106964 562430
rect 107672 555626 107700 568126
rect 110420 566568 110472 566574
rect 110420 566510 110472 566516
rect 108396 565412 108448 565418
rect 108396 565354 108448 565360
rect 108304 565140 108356 565146
rect 108304 565082 108356 565088
rect 107660 555620 107712 555626
rect 107660 555562 107712 555568
rect 108212 555484 108264 555490
rect 108212 555426 108264 555432
rect 107568 552696 107620 552702
rect 107568 552638 107620 552644
rect 106924 550520 106976 550526
rect 106924 550462 106976 550468
rect 106096 550180 106148 550186
rect 106096 550122 106148 550128
rect 106832 550180 106884 550186
rect 106832 550122 106884 550128
rect 106108 547963 106136 550122
rect 106844 547963 106872 550122
rect 107580 547963 107608 552638
rect 108224 547963 108252 555426
rect 108316 550594 108344 565082
rect 108304 550588 108356 550594
rect 108304 550530 108356 550536
rect 108408 550458 108436 565354
rect 109684 565276 109736 565282
rect 109684 565218 109736 565224
rect 109696 557534 109724 565218
rect 109696 557506 109816 557534
rect 109684 550588 109736 550594
rect 109684 550530 109736 550536
rect 108948 550520 109000 550526
rect 108948 550462 109000 550468
rect 108396 550452 108448 550458
rect 108396 550394 108448 550400
rect 108960 547963 108988 550462
rect 109696 547963 109724 550530
rect 109788 549438 109816 557506
rect 110432 552702 110460 566510
rect 110512 565140 110564 565146
rect 110512 565082 110564 565088
rect 110420 552696 110472 552702
rect 110420 552638 110472 552644
rect 109776 549432 109828 549438
rect 109776 549374 109828 549380
rect 110524 548162 110552 565082
rect 110616 554130 110644 568126
rect 112444 565208 112496 565214
rect 112444 565150 112496 565156
rect 111892 562488 111944 562494
rect 111892 562430 111944 562436
rect 110604 554124 110656 554130
rect 110604 554066 110656 554072
rect 111904 552786 111932 562430
rect 112456 552906 112484 565150
rect 113192 557534 113220 568414
rect 114572 568126 114770 568154
rect 117346 568126 117452 568154
rect 114572 562358 114600 568126
rect 115204 565480 115256 565486
rect 115204 565422 115256 565428
rect 114652 565344 114704 565350
rect 114652 565286 114704 565292
rect 114560 562352 114612 562358
rect 114560 562294 114612 562300
rect 113192 557506 113312 557534
rect 112444 552900 112496 552906
rect 112444 552842 112496 552848
rect 111904 552758 112576 552786
rect 111064 552696 111116 552702
rect 111064 552638 111116 552644
rect 110448 548134 110552 548162
rect 110448 547944 110476 548134
rect 111076 547963 111104 552638
rect 111800 550452 111852 550458
rect 111800 550394 111852 550400
rect 111812 547963 111840 550394
rect 112548 547963 112576 552758
rect 113284 547963 113312 557506
rect 114664 550474 114692 565286
rect 115216 550594 115244 565422
rect 117424 565214 117452 568126
rect 120184 568126 120566 568154
rect 117412 565208 117464 565214
rect 117412 565150 117464 565156
rect 120184 564466 120212 568126
rect 120736 565146 120764 630414
rect 120814 606384 120870 606393
rect 120814 606319 120870 606328
rect 120724 565140 120776 565146
rect 120724 565082 120776 565088
rect 116584 564460 116636 564466
rect 116584 564402 116636 564408
rect 120172 564460 120224 564466
rect 120172 564402 120224 564408
rect 116596 552770 116624 564402
rect 118700 562352 118752 562358
rect 118700 562294 118752 562300
rect 118712 557534 118740 562294
rect 120828 558278 120856 606319
rect 120920 568070 120948 633966
rect 122932 633956 122984 633962
rect 122932 633898 122984 633904
rect 140780 633956 140832 633962
rect 140780 633898 140832 633904
rect 121000 633752 121052 633758
rect 121000 633694 121052 633700
rect 120908 568064 120960 568070
rect 120908 568006 120960 568012
rect 121012 568002 121040 633694
rect 122196 633684 122248 633690
rect 122196 633626 122248 633632
rect 121644 633548 121696 633554
rect 121644 633490 121696 633496
rect 121460 630420 121512 630426
rect 121460 630362 121512 630368
rect 121090 591220 121146 591229
rect 121090 591155 121146 591164
rect 121000 567996 121052 568002
rect 121000 567938 121052 567944
rect 120816 558272 120868 558278
rect 120816 558214 120868 558220
rect 118712 557506 119752 557534
rect 116584 552764 116636 552770
rect 116584 552706 116636 552712
rect 115204 550588 115256 550594
rect 115204 550530 115256 550536
rect 116124 550588 116176 550594
rect 116124 550530 116176 550536
rect 114664 550446 115428 550474
rect 114008 550248 114060 550254
rect 114008 550190 114060 550196
rect 114020 547963 114048 550190
rect 114652 549432 114704 549438
rect 114652 549374 114704 549380
rect 114664 547963 114692 549374
rect 115400 547963 115428 550446
rect 116136 547963 116164 550530
rect 116860 549976 116912 549982
rect 116860 549918 116912 549924
rect 116872 547963 116900 549918
rect 117596 549908 117648 549914
rect 117596 549850 117648 549856
rect 118976 549908 119028 549914
rect 118976 549850 119028 549856
rect 117608 547963 117636 549850
rect 118240 549364 118292 549370
rect 118240 549306 118292 549312
rect 118252 547963 118280 549306
rect 118988 547963 119016 549850
rect 119724 547963 119752 557506
rect 121104 557054 121132 591155
rect 121182 578980 121238 578989
rect 121182 578915 121238 578924
rect 121196 562426 121224 578915
rect 121472 576854 121500 630362
rect 121472 576826 121592 576854
rect 121564 570194 121592 576826
rect 121380 570166 121592 570194
rect 121380 568206 121408 570166
rect 121550 570072 121606 570081
rect 121550 570007 121606 570016
rect 121368 568200 121420 568206
rect 121368 568142 121420 568148
rect 121460 568064 121512 568070
rect 121460 568006 121512 568012
rect 121184 562420 121236 562426
rect 121184 562362 121236 562368
rect 121092 557048 121144 557054
rect 121092 556990 121144 556996
rect 121092 556912 121144 556918
rect 121092 556854 121144 556860
rect 120448 551404 120500 551410
rect 120448 551346 120500 551352
rect 120460 547963 120488 551346
rect 121104 547963 121132 556854
rect 121472 552634 121500 568006
rect 121564 567934 121592 570007
rect 121552 567928 121604 567934
rect 121552 567870 121604 567876
rect 121460 552628 121512 552634
rect 121460 552570 121512 552576
rect 121656 550322 121684 633490
rect 121826 621208 121882 621217
rect 121826 621143 121882 621152
rect 121734 615632 121790 615641
rect 121734 615567 121790 615576
rect 121748 554062 121776 615567
rect 121840 559638 121868 621143
rect 121918 608968 121974 608977
rect 121918 608903 121974 608912
rect 121932 561066 121960 608903
rect 122010 594008 122066 594017
rect 122010 593943 122066 593952
rect 122024 566506 122052 593943
rect 122102 588024 122158 588033
rect 122102 587959 122158 587968
rect 122116 566642 122144 587959
rect 122104 566636 122156 566642
rect 122104 566578 122156 566584
rect 122012 566500 122064 566506
rect 122012 566442 122064 566448
rect 121920 561060 121972 561066
rect 121920 561002 121972 561008
rect 121828 559632 121880 559638
rect 121828 559574 121880 559580
rect 121736 554056 121788 554062
rect 121736 553998 121788 554004
rect 121828 552696 121880 552702
rect 121828 552638 121880 552644
rect 121644 550316 121696 550322
rect 121644 550258 121696 550264
rect 121840 547963 121868 552638
rect 122208 550050 122236 633626
rect 122838 628008 122894 628017
rect 122838 627943 122894 627952
rect 122286 572792 122342 572801
rect 122286 572727 122342 572736
rect 122300 568478 122328 572727
rect 122288 568472 122340 568478
rect 122288 568414 122340 568420
rect 122852 560998 122880 627943
rect 122944 568274 122972 633898
rect 124312 633888 124364 633894
rect 124312 633830 124364 633836
rect 124220 630828 124272 630834
rect 124220 630770 124272 630776
rect 123022 625288 123078 625297
rect 123022 625223 123078 625232
rect 122932 568268 122984 568274
rect 122932 568210 122984 568216
rect 123036 562494 123064 625223
rect 123114 612776 123170 612785
rect 123114 612711 123170 612720
rect 123024 562488 123076 562494
rect 123024 562430 123076 562436
rect 122840 560992 122892 560998
rect 122840 560934 122892 560940
rect 122840 559632 122892 559638
rect 122840 559574 122892 559580
rect 122852 552770 122880 559574
rect 123128 559570 123156 612711
rect 123298 603120 123354 603129
rect 123298 603055 123354 603064
rect 123206 600400 123262 600409
rect 123206 600335 123262 600344
rect 123116 559564 123168 559570
rect 123116 559506 123168 559512
rect 122932 558272 122984 558278
rect 122932 558214 122984 558220
rect 122944 552786 122972 558214
rect 123220 557534 123248 600335
rect 123312 558346 123340 603055
rect 124126 596728 124182 596737
rect 124126 596663 124182 596672
rect 124140 596222 124168 596663
rect 124128 596216 124180 596222
rect 124128 596158 124180 596164
rect 123390 584488 123446 584497
rect 123390 584423 123446 584432
rect 123404 563786 123432 584423
rect 123482 581768 123538 581777
rect 123482 581703 123538 581712
rect 123496 576854 123524 581703
rect 123496 576826 123616 576854
rect 123482 575648 123538 575657
rect 123482 575583 123538 575592
rect 123496 567866 123524 575583
rect 123588 568342 123616 576826
rect 123576 568336 123628 568342
rect 123576 568278 123628 568284
rect 123484 567860 123536 567866
rect 123484 567802 123536 567808
rect 123392 563780 123444 563786
rect 123392 563722 123444 563728
rect 123300 558340 123352 558346
rect 123300 558282 123352 558288
rect 123220 557506 123432 557534
rect 122840 552764 122892 552770
rect 122944 552758 123340 552786
rect 122840 552706 122892 552712
rect 122564 552628 122616 552634
rect 122564 552570 122616 552576
rect 122196 550044 122248 550050
rect 122196 549986 122248 549992
rect 122576 547963 122604 552570
rect 123312 547963 123340 552758
rect 123404 551342 123432 557506
rect 124232 552770 124260 630770
rect 124036 552764 124088 552770
rect 124036 552706 124088 552712
rect 124220 552764 124272 552770
rect 124220 552706 124272 552712
rect 123392 551336 123444 551342
rect 123392 551278 123444 551284
rect 124048 547963 124076 552706
rect 124324 550118 124352 633830
rect 124588 633820 124640 633826
rect 124588 633762 124640 633768
rect 124496 633616 124548 633622
rect 124496 633558 124548 633564
rect 124404 630964 124456 630970
rect 124404 630906 124456 630912
rect 124416 550186 124444 630906
rect 124508 568138 124536 633558
rect 124600 568410 124628 633762
rect 133880 633548 133932 633554
rect 133880 633490 133932 633496
rect 124864 631236 124916 631242
rect 124864 631178 124916 631184
rect 124588 568404 124640 568410
rect 124588 568346 124640 568352
rect 124496 568132 124548 568138
rect 124496 568074 124548 568080
rect 124680 551336 124732 551342
rect 124680 551278 124732 551284
rect 124404 550180 124456 550186
rect 124404 550122 124456 550128
rect 124312 550112 124364 550118
rect 124312 550054 124364 550060
rect 124692 547963 124720 551278
rect 124876 549370 124904 631178
rect 125784 630760 125836 630766
rect 125784 630702 125836 630708
rect 125600 585200 125652 585206
rect 125600 585142 125652 585148
rect 125612 555830 125640 585142
rect 125692 566704 125744 566710
rect 125692 566646 125744 566652
rect 125600 555824 125652 555830
rect 125600 555766 125652 555772
rect 125416 552764 125468 552770
rect 125416 552706 125468 552712
rect 124864 549364 124916 549370
rect 124864 549306 124916 549312
rect 125428 547963 125456 552706
rect 125704 550066 125732 566646
rect 125796 550254 125824 630702
rect 132500 615528 132552 615534
rect 132500 615470 132552 615476
rect 129004 597576 129056 597582
rect 129004 597518 129056 597524
rect 126980 563848 127032 563854
rect 126980 563790 127032 563796
rect 126888 555824 126940 555830
rect 126888 555766 126940 555772
rect 125784 550248 125836 550254
rect 125784 550190 125836 550196
rect 125704 550038 126192 550066
rect 126164 547963 126192 550038
rect 126900 547963 126928 555766
rect 126992 552770 127020 563790
rect 129016 557534 129044 597518
rect 130384 582412 130436 582418
rect 130384 582354 130436 582360
rect 129740 565276 129792 565282
rect 129740 565218 129792 565224
rect 128924 557506 129044 557534
rect 127624 554124 127676 554130
rect 127624 554066 127676 554072
rect 126980 552764 127032 552770
rect 126980 552706 127032 552712
rect 127636 547963 127664 554066
rect 128268 552764 128320 552770
rect 128268 552706 128320 552712
rect 128280 547963 128308 552706
rect 128924 549914 128952 557506
rect 129752 552786 129780 565218
rect 130396 557534 130424 582354
rect 131120 558204 131172 558210
rect 131120 558146 131172 558152
rect 131132 557534 131160 558146
rect 130396 557506 130608 557534
rect 131132 557506 131252 557534
rect 129752 552758 130516 552786
rect 129740 552696 129792 552702
rect 129740 552638 129792 552644
rect 129004 549976 129056 549982
rect 129004 549918 129056 549924
rect 128912 549908 128964 549914
rect 128912 549850 128964 549856
rect 129016 547963 129044 549918
rect 129752 547963 129780 552638
rect 130488 547963 130516 552758
rect 130580 551410 130608 557506
rect 130568 551404 130620 551410
rect 130568 551346 130620 551352
rect 131224 547963 131252 557506
rect 132512 552786 132540 615470
rect 132592 565208 132644 565214
rect 132592 565150 132644 565156
rect 132604 557534 132632 565150
rect 132604 557506 133368 557534
rect 132512 552758 132632 552786
rect 131856 549908 131908 549914
rect 131856 549850 131908 549856
rect 131868 547963 131896 549850
rect 132604 547963 132632 552758
rect 133340 547963 133368 557506
rect 133892 557002 133920 633490
rect 136640 630964 136692 630970
rect 136640 630906 136692 630912
rect 133972 565140 134024 565146
rect 133972 565082 134024 565088
rect 133984 557534 134012 565082
rect 136652 557534 136680 630906
rect 140044 630896 140096 630902
rect 140044 630838 140096 630844
rect 139400 579692 139452 579698
rect 139400 579634 139452 579640
rect 138020 561128 138072 561134
rect 138020 561070 138072 561076
rect 138032 557534 138060 561070
rect 139412 557534 139440 579634
rect 133984 557506 134748 557534
rect 136652 557506 137692 557534
rect 138032 557506 138336 557534
rect 139412 557506 139808 557534
rect 133892 556974 134104 557002
rect 134076 547963 134104 556974
rect 134720 547963 134748 557506
rect 137192 556980 137244 556986
rect 137192 556922 137244 556928
rect 135444 551540 135496 551546
rect 135444 551482 135496 551488
rect 135456 547963 135484 551482
rect 136180 550588 136232 550594
rect 136180 550530 136232 550536
rect 136192 547963 136220 550530
rect 136916 550044 136968 550050
rect 136916 549986 136968 549992
rect 136928 547963 136956 549986
rect 137204 549982 137232 556922
rect 137192 549976 137244 549982
rect 137192 549918 137244 549924
rect 137664 547963 137692 557506
rect 138308 547963 138336 557506
rect 139032 550112 139084 550118
rect 139032 550054 139084 550060
rect 139044 547963 139072 550054
rect 139780 547963 139808 557506
rect 140056 550594 140084 630838
rect 140504 554056 140556 554062
rect 140504 553998 140556 554004
rect 140044 550588 140096 550594
rect 140044 550530 140096 550536
rect 140516 547963 140544 553998
rect 140792 552770 140820 633898
rect 142160 633752 142212 633758
rect 142160 633694 142212 633700
rect 140872 619676 140924 619682
rect 140872 619618 140924 619624
rect 140884 557534 140912 619618
rect 140884 557506 141280 557534
rect 140780 552764 140832 552770
rect 140780 552706 140832 552712
rect 141252 547963 141280 557506
rect 142172 552770 142200 633694
rect 144184 631100 144236 631106
rect 144184 631042 144236 631048
rect 143540 565480 143592 565486
rect 143540 565422 143592 565428
rect 142620 555620 142672 555626
rect 142620 555562 142672 555568
rect 141884 552764 141936 552770
rect 141884 552706 141936 552712
rect 142160 552764 142212 552770
rect 142160 552706 142212 552712
rect 141896 547963 141924 552706
rect 142632 547963 142660 555562
rect 143552 552770 143580 565422
rect 143356 552764 143408 552770
rect 143356 552706 143408 552712
rect 143540 552764 143592 552770
rect 143540 552706 143592 552712
rect 143368 547963 143396 552706
rect 144092 550384 144144 550390
rect 144092 550326 144144 550332
rect 144104 547963 144132 550326
rect 144196 549914 144224 631042
rect 144276 627972 144328 627978
rect 144276 627914 144328 627920
rect 144288 551546 144316 627914
rect 144932 552770 144960 634102
rect 145012 634092 145064 634098
rect 145012 634034 145064 634040
rect 145024 557534 145052 634034
rect 147496 633616 147548 633622
rect 147496 633558 147548 633564
rect 147404 633480 147456 633486
rect 147404 633422 147456 633428
rect 146116 631304 146168 631310
rect 146116 631246 146168 631252
rect 145564 596216 145616 596222
rect 145564 596158 145616 596164
rect 145576 568478 145604 596158
rect 145564 568472 145616 568478
rect 145564 568414 145616 568420
rect 145024 557506 145512 557534
rect 144736 552764 144788 552770
rect 144736 552706 144788 552712
rect 144920 552764 144972 552770
rect 144920 552706 144972 552712
rect 144276 551540 144328 551546
rect 144276 551482 144328 551488
rect 144184 549908 144236 549914
rect 144184 549850 144236 549856
rect 144748 547963 144776 552706
rect 145484 547963 145512 557506
rect 146128 550254 146156 631246
rect 146208 630692 146260 630698
rect 146208 630634 146260 630640
rect 146220 604217 146248 630634
rect 146298 628688 146354 628697
rect 146298 628623 146354 628632
rect 146312 627978 146340 628623
rect 146300 627972 146352 627978
rect 146300 627914 146352 627920
rect 147310 622432 147366 622441
rect 147310 622367 147366 622376
rect 146298 619712 146354 619721
rect 146298 619647 146300 619656
rect 146352 619647 146354 619656
rect 146300 619618 146352 619624
rect 146298 616312 146354 616321
rect 146298 616247 146354 616256
rect 146312 615534 146340 616247
rect 146300 615528 146352 615534
rect 146300 615470 146352 615476
rect 146850 613592 146906 613601
rect 146850 613527 146906 613536
rect 146206 604208 146262 604217
rect 146206 604143 146262 604152
rect 146298 597952 146354 597961
rect 146298 597887 146354 597896
rect 146312 597582 146340 597887
rect 146300 597576 146352 597582
rect 146300 597518 146352 597524
rect 146298 585712 146354 585721
rect 146298 585647 146354 585656
rect 146312 585206 146340 585647
rect 146300 585200 146352 585206
rect 146300 585142 146352 585148
rect 146298 582992 146354 583001
rect 146298 582927 146354 582936
rect 146312 582418 146340 582927
rect 146300 582412 146352 582418
rect 146300 582354 146352 582360
rect 146298 579728 146354 579737
rect 146298 579663 146300 579672
rect 146352 579663 146354 579672
rect 146300 579634 146352 579640
rect 146864 563786 146892 613527
rect 147126 595232 147182 595241
rect 147126 595167 147182 595176
rect 147034 576872 147090 576881
rect 147034 576807 147090 576816
rect 146852 563780 146904 563786
rect 146852 563722 146904 563728
rect 147048 561066 147076 576807
rect 147140 568410 147168 595167
rect 147218 589112 147274 589121
rect 147218 589047 147274 589056
rect 147128 568404 147180 568410
rect 147128 568346 147180 568352
rect 147036 561060 147088 561066
rect 147036 561002 147088 561008
rect 147232 556850 147260 589047
rect 147324 560998 147352 622367
rect 147416 568002 147444 633422
rect 147508 568138 147536 633558
rect 147600 607617 147628 683130
rect 299492 641034 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 305644 700460 305696 700466
rect 305644 700402 305696 700408
rect 299480 641028 299532 641034
rect 299480 640970 299532 640976
rect 236644 634228 236696 634234
rect 236644 634170 236696 634176
rect 156604 634092 156656 634098
rect 156604 634034 156656 634040
rect 207664 634092 207716 634098
rect 207664 634034 207716 634040
rect 148876 634024 148928 634030
rect 148876 633966 148928 633972
rect 148784 633888 148836 633894
rect 148784 633830 148836 633836
rect 148324 630760 148376 630766
rect 148324 630702 148376 630708
rect 147586 607608 147642 607617
rect 147586 607543 147642 607552
rect 148230 570752 148286 570761
rect 148230 570687 148286 570696
rect 147496 568132 147548 568138
rect 147496 568074 147548 568080
rect 147404 567996 147456 568002
rect 147404 567938 147456 567944
rect 148244 561202 148272 570687
rect 148232 561196 148284 561202
rect 148232 561138 148284 561144
rect 147312 560992 147364 560998
rect 147312 560934 147364 560940
rect 147220 556844 147272 556850
rect 147220 556786 147272 556792
rect 146300 552832 146352 552838
rect 146300 552774 146352 552780
rect 146208 552764 146260 552770
rect 146208 552706 146260 552712
rect 146116 550248 146168 550254
rect 146116 550190 146168 550196
rect 146220 547963 146248 552706
rect 146312 550390 146340 552774
rect 147680 551540 147732 551546
rect 147680 551482 147732 551488
rect 146944 550588 146996 550594
rect 146944 550530 146996 550536
rect 146300 550384 146352 550390
rect 146300 550326 146352 550332
rect 146956 547963 146984 550530
rect 147692 547963 147720 551482
rect 148336 550594 148364 630702
rect 148690 625832 148746 625841
rect 148690 625767 148746 625776
rect 148506 610192 148562 610201
rect 148506 610127 148562 610136
rect 148414 591832 148470 591841
rect 148414 591767 148470 591776
rect 148428 552022 148456 591767
rect 148520 566506 148548 610127
rect 148598 601352 148654 601361
rect 148598 601287 148654 601296
rect 148508 566500 148560 566506
rect 148508 566442 148560 566448
rect 148508 552764 148560 552770
rect 148508 552706 148560 552712
rect 148416 552016 148468 552022
rect 148416 551958 148468 551964
rect 148324 550588 148376 550594
rect 148324 550530 148376 550536
rect 148520 548162 148548 552706
rect 148612 551954 148640 601287
rect 148704 565894 148732 625767
rect 148796 567934 148824 633830
rect 148784 567928 148836 567934
rect 148784 567870 148836 567876
rect 148888 567866 148916 633966
rect 149796 633820 149848 633826
rect 149796 633762 149848 633768
rect 149704 633480 149756 633486
rect 149704 633422 149756 633428
rect 148968 631168 149020 631174
rect 148968 631110 149020 631116
rect 148876 567860 148928 567866
rect 148876 567802 148928 567808
rect 148692 565888 148744 565894
rect 148692 565830 148744 565836
rect 148600 551948 148652 551954
rect 148600 551890 148652 551896
rect 148980 549914 149008 631110
rect 149058 573472 149114 573481
rect 149058 573407 149114 573416
rect 149072 559570 149100 573407
rect 149716 568206 149744 633422
rect 149704 568200 149756 568206
rect 149704 568142 149756 568148
rect 149808 567254 149836 633762
rect 156616 633690 156644 634034
rect 172888 634024 172940 634030
rect 172888 633966 172940 633972
rect 167092 633956 167144 633962
rect 167092 633898 167144 633904
rect 156604 633684 156656 633690
rect 156604 633626 156656 633632
rect 149980 633548 150032 633554
rect 149980 633490 150032 633496
rect 149888 631032 149940 631038
rect 149888 630974 149940 630980
rect 149992 630986 150020 633490
rect 164516 633480 164568 633486
rect 164516 633422 164568 633428
rect 155500 631304 155552 631310
rect 155500 631246 155552 631252
rect 155512 630986 155540 631246
rect 158720 631168 158772 631174
rect 158720 631110 158772 631116
rect 158732 630986 158760 631110
rect 161480 631100 161532 631106
rect 161480 631042 161532 631048
rect 161492 630986 161520 631042
rect 164528 630986 164556 633422
rect 167104 630986 167132 633898
rect 170312 631032 170364 631038
rect 149796 567248 149848 567254
rect 149796 567190 149848 567196
rect 149060 559564 149112 559570
rect 149060 559506 149112 559512
rect 149060 552016 149112 552022
rect 149060 551958 149112 551964
rect 148968 549908 149020 549914
rect 148968 549850 149020 549856
rect 148352 548134 148548 548162
rect 148352 547944 148380 548134
rect 149072 547963 149100 551958
rect 149796 551948 149848 551954
rect 149796 551890 149848 551896
rect 149808 547963 149836 551890
rect 149900 550594 149928 630974
rect 149992 630958 150052 630986
rect 155512 630958 155848 630986
rect 158732 630958 159068 630986
rect 161492 630958 161644 630986
rect 164528 630958 164864 630986
rect 167104 630958 167440 630986
rect 172900 630986 172928 633966
rect 176108 633888 176160 633894
rect 176108 633830 176160 633836
rect 176120 630986 176148 633830
rect 190552 633820 190604 633826
rect 190552 633762 190604 633768
rect 184480 633752 184532 633758
rect 184480 633694 184532 633700
rect 184492 630986 184520 633694
rect 187700 631236 187752 631242
rect 187700 631178 187752 631184
rect 187712 630986 187740 631178
rect 190564 630986 190592 633762
rect 196072 633684 196124 633690
rect 196072 633626 196124 633632
rect 196084 630986 196112 633626
rect 199292 633616 199344 633622
rect 199292 633558 199344 633564
rect 199304 630986 199332 633558
rect 201868 633548 201920 633554
rect 201868 633490 201920 633496
rect 205548 633548 205600 633554
rect 205548 633490 205600 633496
rect 201880 630986 201908 633490
rect 205560 630986 205588 633490
rect 170364 630980 170660 630986
rect 170312 630974 170660 630980
rect 170324 630958 170660 630974
rect 172900 630958 173236 630986
rect 176120 630958 176456 630986
rect 178696 630970 179032 630986
rect 178684 630964 179032 630970
rect 178736 630958 179032 630964
rect 184492 630958 184828 630986
rect 187712 630958 188048 630986
rect 190564 630958 190624 630986
rect 196084 630958 196420 630986
rect 199304 630958 199640 630986
rect 201880 630958 202216 630986
rect 205436 630958 205588 630986
rect 207676 630986 207704 634034
rect 226340 634024 226392 634030
rect 226340 633966 226392 633972
rect 214012 633956 214064 633962
rect 214012 633898 214064 633904
rect 213920 633684 213972 633690
rect 213920 633626 213972 633632
rect 212632 633548 212684 633554
rect 212632 633490 212684 633496
rect 207676 630958 208012 630986
rect 178684 630906 178736 630912
rect 193496 630896 193548 630902
rect 182100 630834 182252 630850
rect 193548 630844 193844 630850
rect 193496 630838 193844 630844
rect 182088 630828 182252 630834
rect 182140 630822 182252 630828
rect 193508 630822 193844 630838
rect 182088 630770 182140 630776
rect 153108 630760 153160 630766
rect 153160 630708 153272 630714
rect 153108 630702 153272 630708
rect 153120 630686 153272 630702
rect 210588 630414 210740 630442
rect 151084 568404 151136 568410
rect 151084 568346 151136 568352
rect 150052 568126 150388 568154
rect 150360 564602 150388 568126
rect 150532 565888 150584 565894
rect 150532 565830 150584 565836
rect 150348 564596 150400 564602
rect 150348 564538 150400 564544
rect 149888 550588 149940 550594
rect 149888 550530 149940 550536
rect 150544 547963 150572 565830
rect 151096 550390 151124 568346
rect 154764 568200 154816 568206
rect 151924 568126 152628 568154
rect 204904 568200 204956 568206
rect 154764 568142 154816 568148
rect 151820 567248 151872 567254
rect 151820 567190 151872 567196
rect 151176 564596 151228 564602
rect 151176 564538 151228 564544
rect 151188 554198 151216 564538
rect 151176 554192 151228 554198
rect 151176 554134 151228 554140
rect 151832 552786 151860 567190
rect 151924 557534 151952 568126
rect 154672 565412 154724 565418
rect 154672 565354 154724 565360
rect 151924 557506 152044 557534
rect 151832 552758 151952 552786
rect 151268 550588 151320 550594
rect 151268 550530 151320 550536
rect 151084 550384 151136 550390
rect 151084 550326 151136 550332
rect 151280 547963 151308 550530
rect 151924 547963 151952 552758
rect 152016 550186 152044 557506
rect 154684 552786 154712 565354
rect 154776 557534 154804 568142
rect 154868 568126 155204 568154
rect 156052 568132 156104 568138
rect 154868 562358 154896 568126
rect 156052 568074 156104 568080
rect 157444 568126 158424 568154
rect 160112 568126 161000 568154
rect 163884 568126 164220 568154
rect 164424 568132 164476 568138
rect 154856 562352 154908 562358
rect 154856 562294 154908 562300
rect 156064 557534 156092 568074
rect 157340 567996 157392 568002
rect 157340 567938 157392 567944
rect 156604 566772 156656 566778
rect 156604 566714 156656 566720
rect 154776 557506 155540 557534
rect 156064 557506 156276 557534
rect 154684 552758 154896 552786
rect 152648 551472 152700 551478
rect 152648 551414 152700 551420
rect 152004 550180 152056 550186
rect 152004 550122 152056 550128
rect 152660 547963 152688 551414
rect 153384 550384 153436 550390
rect 153384 550326 153436 550332
rect 153396 547963 153424 550326
rect 154120 549976 154172 549982
rect 154120 549918 154172 549924
rect 154132 547963 154160 549918
rect 154868 547963 154896 552758
rect 155512 547963 155540 557506
rect 156248 547963 156276 557506
rect 156616 550050 156644 566714
rect 157352 552786 157380 567938
rect 157444 553874 157472 568126
rect 158720 565344 158772 565350
rect 158720 565286 158772 565292
rect 157524 562556 157576 562562
rect 157524 562498 157576 562504
rect 157536 557534 157564 562498
rect 157536 557506 158392 557534
rect 157444 553846 157840 553874
rect 157352 552758 157748 552786
rect 156972 550248 157024 550254
rect 156972 550190 157024 550196
rect 156604 550044 156656 550050
rect 156604 549986 156656 549992
rect 156984 547963 157012 550190
rect 157720 547963 157748 552758
rect 157812 550322 157840 553846
rect 157800 550316 157852 550322
rect 157800 550258 157852 550264
rect 158364 547963 158392 557506
rect 158732 552702 158760 565286
rect 158812 561196 158864 561202
rect 158812 561138 158864 561144
rect 158824 557534 158852 561138
rect 158824 557506 159128 557534
rect 158720 552696 158772 552702
rect 158720 552638 158772 552644
rect 159100 547963 159128 557506
rect 159824 552696 159876 552702
rect 159824 552638 159876 552644
rect 159836 547963 159864 552638
rect 160112 550050 160140 568126
rect 161480 567928 161532 567934
rect 161480 567870 161532 567876
rect 160192 566500 160244 566506
rect 160192 566442 160244 566448
rect 160204 552786 160232 566442
rect 160284 559564 160336 559570
rect 160284 559506 160336 559512
rect 160296 557534 160324 559506
rect 160296 557506 161336 557534
rect 160204 552758 160600 552786
rect 160100 550044 160152 550050
rect 160100 549986 160152 549992
rect 160572 547963 160600 552758
rect 161308 547963 161336 557506
rect 161492 552786 161520 567870
rect 161572 565616 161624 565622
rect 161572 565558 161624 565564
rect 161584 557534 161612 565558
rect 163044 565548 163096 565554
rect 163044 565490 163096 565496
rect 163056 557534 163084 565490
rect 163884 565282 163912 568126
rect 164424 568074 164476 568080
rect 166460 568126 166796 568154
rect 169772 568126 170016 568154
rect 172532 568126 172592 568154
rect 175292 568126 175812 568154
rect 178052 568126 178388 568154
rect 181272 568126 181608 568154
rect 183848 568126 184184 568154
rect 187068 568126 187404 568154
rect 189644 568126 189980 568154
rect 192864 568126 193200 568154
rect 195440 568126 195776 568154
rect 198752 568126 198996 568154
rect 201512 568126 201572 568154
rect 204456 568126 204792 568154
rect 204904 568142 204956 568148
rect 164332 567860 164384 567866
rect 164332 567802 164384 567808
rect 163872 565276 163924 565282
rect 163872 565218 163924 565224
rect 161584 557506 162716 557534
rect 163056 557506 164188 557534
rect 161492 552758 161980 552786
rect 161952 547963 161980 552758
rect 162688 547963 162716 557506
rect 163412 554192 163464 554198
rect 163412 554134 163464 554140
rect 163424 547963 163452 554134
rect 164160 547963 164188 557506
rect 164344 552786 164372 567802
rect 164436 557534 164464 568074
rect 166460 565486 166488 568126
rect 166448 565480 166500 565486
rect 166448 565422 166500 565428
rect 165620 563780 165672 563786
rect 165620 563722 165672 563728
rect 165632 557534 165660 563722
rect 168380 561060 168432 561066
rect 168380 561002 168432 561008
rect 168392 557534 168420 561002
rect 164436 557506 165568 557534
rect 165632 557506 166304 557534
rect 168392 557506 169156 557534
rect 164344 552758 164924 552786
rect 164896 547963 164924 552758
rect 165540 547963 165568 557506
rect 166276 547963 166304 557506
rect 168380 554260 168432 554266
rect 168380 554202 168432 554208
rect 167000 550316 167052 550322
rect 167000 550258 167052 550264
rect 167012 547963 167040 550258
rect 167736 550180 167788 550186
rect 167736 550122 167788 550128
rect 167748 547963 167776 550122
rect 168392 547963 168420 554202
rect 169128 547963 169156 557506
rect 169772 549846 169800 568126
rect 172532 552770 172560 568126
rect 173900 565480 173952 565486
rect 173900 565422 173952 565428
rect 173912 557534 173940 565422
rect 173912 557506 174216 557534
rect 173808 552968 173860 552974
rect 173808 552910 173860 552916
rect 172520 552764 172572 552770
rect 172520 552706 172572 552712
rect 173820 550458 173848 552910
rect 171324 550452 171376 550458
rect 171324 550394 171376 550400
rect 173808 550452 173860 550458
rect 173808 550394 173860 550400
rect 169852 550248 169904 550254
rect 169852 550190 169904 550196
rect 169760 549840 169812 549846
rect 169760 549782 169812 549788
rect 169864 547963 169892 550190
rect 170588 550180 170640 550186
rect 170588 550122 170640 550128
rect 170600 547963 170628 550122
rect 171336 547963 171364 550394
rect 172704 550044 172756 550050
rect 172704 549986 172756 549992
rect 171968 549908 172020 549914
rect 171968 549850 172020 549856
rect 171980 547963 172008 549850
rect 172716 547963 172744 549986
rect 173440 549840 173492 549846
rect 173440 549782 173492 549788
rect 173452 547963 173480 549782
rect 174188 547963 174216 557506
rect 174912 556844 174964 556850
rect 174912 556786 174964 556792
rect 174924 547963 174952 556786
rect 175292 550254 175320 568126
rect 178052 565622 178080 568126
rect 179420 567860 179472 567866
rect 179420 567802 179472 567808
rect 178040 565616 178092 565622
rect 178040 565558 178092 565564
rect 176660 561196 176712 561202
rect 176660 561138 176712 561144
rect 175372 560992 175424 560998
rect 175372 560934 175424 560940
rect 175384 557534 175412 560934
rect 175384 557506 175596 557534
rect 175280 550248 175332 550254
rect 175280 550190 175332 550196
rect 175568 547963 175596 557506
rect 176672 552786 176700 561138
rect 176752 559768 176804 559774
rect 176752 559710 176804 559716
rect 176764 557534 176792 559710
rect 178040 558408 178092 558414
rect 178040 558350 178092 558356
rect 178052 557534 178080 558350
rect 176764 557506 177804 557534
rect 178052 557506 178540 557534
rect 176672 552758 177068 552786
rect 176292 549908 176344 549914
rect 176292 549850 176344 549856
rect 176304 547963 176332 549850
rect 177040 547963 177068 552758
rect 177776 547963 177804 557506
rect 178512 547963 178540 557506
rect 179144 556844 179196 556850
rect 179144 556786 179196 556792
rect 179156 547963 179184 556786
rect 179432 552770 179460 567802
rect 180984 566568 181036 566574
rect 180984 566510 181036 566516
rect 179512 566500 179564 566506
rect 179512 566442 179564 566448
rect 179524 557534 179552 566442
rect 180892 563780 180944 563786
rect 180892 563722 180944 563728
rect 179524 557506 179920 557534
rect 179420 552764 179472 552770
rect 179420 552706 179472 552712
rect 179892 547963 179920 557506
rect 180904 552770 180932 563722
rect 180996 557534 181024 566510
rect 181272 565418 181300 568126
rect 183652 567928 183704 567934
rect 183652 567870 183704 567876
rect 181260 565412 181312 565418
rect 181260 565354 181312 565360
rect 182180 560992 182232 560998
rect 182180 560934 182232 560940
rect 182192 557534 182220 560934
rect 180996 557506 181392 557534
rect 182192 557506 182772 557534
rect 180616 552764 180668 552770
rect 180616 552706 180668 552712
rect 180892 552764 180944 552770
rect 180892 552706 180944 552712
rect 180628 547963 180656 552706
rect 181364 547963 181392 557506
rect 181996 552764 182048 552770
rect 181996 552706 182048 552712
rect 182008 547963 182036 552706
rect 182744 547963 182772 557506
rect 183664 552752 183692 567870
rect 183848 565554 183876 568126
rect 183836 565548 183888 565554
rect 183836 565490 183888 565496
rect 184204 565276 184256 565282
rect 184204 565218 184256 565224
rect 184216 557534 184244 565218
rect 187068 565214 187096 568126
rect 189644 565486 189672 568126
rect 189632 565480 189684 565486
rect 189632 565422 189684 565428
rect 187792 565412 187844 565418
rect 187792 565354 187844 565360
rect 187056 565208 187108 565214
rect 187056 565150 187108 565156
rect 184940 562420 184992 562426
rect 184940 562362 184992 562368
rect 184952 557534 184980 562362
rect 186320 562352 186372 562358
rect 186320 562294 186372 562300
rect 184216 557506 184336 557534
rect 184952 557506 185624 557534
rect 183664 552724 184244 552752
rect 183468 550044 183520 550050
rect 183468 549986 183520 549992
rect 183480 547963 183508 549986
rect 184216 547963 184244 552724
rect 184308 550118 184336 557506
rect 184940 554192 184992 554198
rect 184940 554134 184992 554140
rect 184296 550112 184348 550118
rect 184296 550054 184348 550060
rect 184952 547963 184980 554134
rect 185596 547963 185624 557506
rect 186332 547963 186360 562294
rect 187700 561060 187752 561066
rect 187700 561002 187752 561008
rect 187712 557534 187740 561002
rect 187804 558210 187832 565354
rect 192864 565350 192892 568126
rect 194784 567996 194836 568002
rect 194784 567938 194836 567944
rect 192852 565344 192904 565350
rect 192852 565286 192904 565292
rect 191104 564460 191156 564466
rect 191104 564402 191156 564408
rect 190460 559700 190512 559706
rect 190460 559642 190512 559648
rect 187792 558204 187844 558210
rect 187792 558146 187844 558152
rect 187712 557506 187832 557534
rect 187056 555484 187108 555490
rect 187056 555426 187108 555432
rect 187068 547963 187096 555426
rect 187804 547963 187832 557506
rect 189908 557048 189960 557054
rect 189908 556990 189960 556996
rect 189172 555552 189224 555558
rect 189172 555494 189224 555500
rect 188528 551404 188580 551410
rect 188528 551346 188580 551352
rect 188540 547963 188568 551346
rect 189184 547963 189212 555494
rect 189920 547963 189948 556990
rect 190472 552770 190500 559642
rect 190552 558476 190604 558482
rect 190552 558418 190604 558424
rect 190564 557534 190592 558418
rect 190564 557506 190684 557534
rect 190460 552764 190512 552770
rect 190460 552706 190512 552712
rect 190656 547963 190684 557506
rect 191116 551546 191144 564402
rect 191840 563916 191892 563922
rect 191840 563858 191892 563864
rect 191852 552786 191880 563858
rect 191932 562488 191984 562494
rect 191932 562430 191984 562436
rect 191944 557534 191972 562430
rect 194796 557534 194824 567938
rect 195244 565208 195296 565214
rect 195244 565150 195296 565156
rect 191944 557506 192800 557534
rect 194796 557506 195008 557534
rect 191380 552764 191432 552770
rect 191852 552758 192156 552786
rect 191380 552706 191432 552712
rect 191104 551540 191156 551546
rect 191104 551482 191156 551488
rect 191392 547963 191420 552706
rect 192128 547963 192156 552758
rect 192772 547963 192800 557506
rect 193496 554396 193548 554402
rect 193496 554338 193548 554344
rect 193508 547963 193536 554338
rect 194232 550112 194284 550118
rect 194232 550054 194284 550060
rect 194244 547963 194272 550054
rect 194980 547963 195008 557506
rect 195256 550186 195284 565150
rect 195440 564466 195468 568126
rect 198752 565418 198780 568126
rect 200120 566636 200172 566642
rect 200120 566578 200172 566584
rect 198740 565412 198792 565418
rect 198740 565354 198792 565360
rect 196624 565344 196676 565350
rect 196624 565286 196676 565292
rect 195428 564460 195480 564466
rect 195428 564402 195480 564408
rect 195980 559564 196032 559570
rect 195980 559506 196032 559512
rect 195992 552770 196020 559506
rect 196072 558204 196124 558210
rect 196072 558146 196124 558152
rect 196084 557534 196112 558146
rect 196084 557506 196388 557534
rect 195980 552764 196032 552770
rect 195980 552706 196032 552712
rect 195612 550248 195664 550254
rect 195612 550190 195664 550196
rect 195244 550180 195296 550186
rect 195244 550122 195296 550128
rect 195624 547963 195652 550190
rect 196360 547963 196388 557506
rect 196636 554062 196664 565286
rect 198004 564460 198056 564466
rect 198004 564402 198056 564408
rect 198016 556918 198044 564402
rect 198740 561264 198792 561270
rect 198740 561206 198792 561212
rect 198004 556912 198056 556918
rect 198004 556854 198056 556860
rect 197820 555688 197872 555694
rect 197820 555630 197872 555636
rect 196624 554056 196676 554062
rect 196624 553998 196676 554004
rect 197084 552764 197136 552770
rect 197084 552706 197136 552712
rect 197096 547963 197124 552706
rect 197832 547963 197860 555630
rect 198556 554056 198608 554062
rect 198556 553998 198608 554004
rect 198568 547963 198596 553998
rect 198752 552770 198780 561206
rect 199200 557116 199252 557122
rect 199200 557058 199252 557064
rect 198740 552764 198792 552770
rect 198740 552706 198792 552712
rect 199212 547963 199240 557058
rect 199936 552764 199988 552770
rect 200132 552752 200160 566578
rect 201512 564466 201540 568126
rect 204456 564466 204484 568126
rect 201500 564460 201552 564466
rect 201500 564402 201552 564408
rect 202144 564460 202196 564466
rect 202144 564402 202196 564408
rect 204444 564460 204496 564466
rect 204444 564402 204496 564408
rect 200212 563984 200264 563990
rect 200212 563926 200264 563932
rect 200224 553110 200252 563926
rect 201500 559836 201552 559842
rect 201500 559778 201552 559784
rect 200212 553104 200264 553110
rect 200212 553046 200264 553052
rect 201408 553104 201460 553110
rect 201408 553046 201460 553052
rect 200132 552724 200712 552752
rect 199936 552706 199988 552712
rect 199948 547963 199976 552706
rect 200684 547963 200712 552724
rect 201420 547963 201448 553046
rect 201512 552770 201540 559778
rect 202156 554130 202184 564402
rect 204260 562624 204312 562630
rect 204260 562566 204312 562572
rect 204272 557534 204300 562566
rect 204272 557506 204852 557534
rect 202236 556912 202288 556918
rect 202236 556854 202288 556860
rect 202144 554124 202196 554130
rect 202144 554066 202196 554072
rect 201500 552764 201552 552770
rect 201500 552706 201552 552712
rect 202248 548162 202276 556854
rect 202788 552764 202840 552770
rect 202788 552706 202840 552712
rect 202172 548134 202276 548162
rect 202172 547944 202200 548134
rect 202800 547963 202828 552706
rect 204260 550384 204312 550390
rect 204260 550326 204312 550332
rect 203524 550316 203576 550322
rect 203524 550258 203576 550264
rect 203536 547963 203564 550258
rect 204272 547963 204300 550326
rect 204824 549794 204852 557506
rect 204916 549982 204944 568142
rect 207032 568126 207368 568154
rect 210252 568126 210588 568154
rect 207032 565146 207060 568126
rect 210252 565350 210280 568126
rect 210240 565344 210292 565350
rect 210240 565286 210292 565292
rect 207020 565140 207072 565146
rect 207020 565082 207072 565088
rect 205640 558340 205692 558346
rect 205640 558282 205692 558288
rect 204904 549976 204956 549982
rect 204904 549918 204956 549924
rect 204824 549766 205036 549794
rect 205008 547963 205036 549766
rect 205652 547963 205680 558282
rect 206376 554328 206428 554334
rect 206376 554270 206428 554276
rect 206388 547963 206416 554270
rect 210712 554266 210740 630414
rect 211250 628008 211306 628017
rect 211250 627943 211306 627952
rect 211158 615632 211214 615641
rect 211158 615567 211214 615576
rect 210790 575648 210846 575657
rect 210790 575583 210846 575592
rect 210700 554260 210752 554266
rect 210700 554202 210752 554208
rect 210804 553042 210832 575583
rect 210882 570344 210938 570353
rect 210882 570279 210938 570288
rect 210792 553036 210844 553042
rect 210792 552978 210844 552984
rect 210700 552628 210752 552634
rect 210700 552570 210752 552576
rect 207112 551676 207164 551682
rect 207112 551618 207164 551624
rect 207124 547963 207152 551618
rect 207848 551608 207900 551614
rect 207848 551550 207900 551556
rect 207860 547963 207888 551550
rect 208584 551540 208636 551546
rect 208584 551482 208636 551488
rect 208596 547963 208624 551482
rect 209228 550452 209280 550458
rect 209228 550394 209280 550400
rect 209240 547963 209268 550394
rect 209964 550180 210016 550186
rect 209964 550122 210016 550128
rect 209976 547963 210004 550122
rect 210712 547963 210740 552570
rect 210896 551342 210924 570279
rect 211172 552906 211200 615567
rect 211264 568070 211292 627943
rect 211434 618488 211490 618497
rect 211434 618423 211490 618432
rect 211342 612776 211398 612785
rect 211342 612711 211398 612720
rect 211252 568064 211304 568070
rect 211252 568006 211304 568012
rect 211356 559638 211384 612711
rect 211448 566710 211476 618423
rect 211618 606384 211674 606393
rect 211618 606319 211674 606328
rect 211526 600400 211582 600409
rect 211526 600335 211582 600344
rect 211436 566704 211488 566710
rect 211436 566646 211488 566652
rect 211344 559632 211396 559638
rect 211344 559574 211396 559580
rect 211160 552900 211212 552906
rect 211160 552842 211212 552848
rect 211436 552016 211488 552022
rect 211436 551958 211488 551964
rect 210884 551336 210936 551342
rect 210884 551278 210936 551284
rect 211448 547963 211476 551958
rect 211540 551478 211568 600335
rect 211632 561134 211660 606319
rect 211710 594008 211766 594017
rect 211710 593943 211766 593952
rect 211620 561128 211672 561134
rect 211620 561070 211672 561076
rect 211724 558278 211752 593943
rect 211802 584488 211858 584497
rect 211802 584423 211858 584432
rect 211816 563854 211844 584423
rect 212538 581768 212594 581777
rect 212538 581703 212594 581712
rect 211804 563848 211856 563854
rect 211804 563790 211856 563796
rect 212552 562562 212580 581703
rect 212644 568138 212672 633490
rect 212722 625288 212778 625297
rect 212722 625223 212778 625232
rect 212632 568132 212684 568138
rect 212632 568074 212684 568080
rect 212736 565214 212764 625223
rect 213274 621208 213330 621217
rect 213274 621143 213330 621152
rect 212814 608968 212870 608977
rect 212814 608903 212870 608912
rect 212724 565208 212776 565214
rect 212724 565150 212776 565156
rect 212540 562556 212592 562562
rect 212540 562498 212592 562504
rect 211712 558272 211764 558278
rect 211712 558214 211764 558220
rect 212828 556986 212856 608903
rect 212906 603120 212962 603129
rect 212906 603055 212962 603064
rect 212920 568206 212948 603055
rect 213090 590744 213146 590753
rect 213090 590679 213146 590688
rect 212998 588024 213054 588033
rect 212998 587959 213054 587968
rect 212908 568200 212960 568206
rect 212908 568142 212960 568148
rect 212816 556980 212868 556986
rect 212816 556922 212868 556928
rect 213012 555626 213040 587959
rect 213104 565282 213132 590679
rect 213182 578368 213238 578377
rect 213182 578303 213238 578312
rect 213196 566778 213224 578303
rect 213184 566772 213236 566778
rect 213184 566714 213236 566720
rect 213092 565276 213144 565282
rect 213092 565218 213144 565224
rect 213000 555620 213052 555626
rect 213000 555562 213052 555568
rect 213288 552838 213316 621143
rect 213366 572792 213422 572801
rect 213366 572727 213422 572736
rect 213380 552974 213408 572727
rect 213552 553036 213604 553042
rect 213552 552978 213604 552984
rect 213368 552968 213420 552974
rect 213368 552910 213420 552916
rect 213276 552832 213328 552838
rect 213276 552774 213328 552780
rect 212172 552696 212224 552702
rect 212172 552638 212224 552644
rect 211528 551472 211580 551478
rect 211528 551414 211580 551420
rect 212184 547963 212212 552638
rect 212816 549976 212868 549982
rect 212816 549918 212868 549924
rect 212828 547963 212856 549918
rect 213564 547963 213592 552978
rect 213932 552770 213960 633626
rect 214024 557534 214052 633898
rect 223580 633004 223632 633010
rect 223580 632946 223632 632952
rect 222200 632936 222252 632942
rect 222200 632878 222252 632884
rect 217324 631032 217376 631038
rect 217324 630974 217376 630980
rect 214564 630964 214616 630970
rect 214564 630906 214616 630912
rect 214102 596728 214158 596737
rect 214102 596663 214158 596672
rect 214116 568478 214144 596663
rect 214104 568472 214156 568478
rect 214104 568414 214156 568420
rect 214024 557506 214328 557534
rect 213920 552764 213972 552770
rect 213920 552706 213972 552712
rect 214300 547963 214328 557506
rect 214576 550254 214604 630906
rect 215944 630760 215996 630766
rect 215944 630702 215996 630708
rect 215300 629944 215352 629950
rect 215300 629886 215352 629892
rect 214656 594856 214708 594862
rect 214656 594798 214708 594804
rect 214668 552022 214696 594798
rect 215312 552786 215340 629886
rect 215392 563848 215444 563854
rect 215392 563790 215444 563796
rect 215404 557534 215432 563790
rect 215404 557506 215892 557534
rect 215024 552764 215076 552770
rect 215312 552758 215800 552786
rect 215024 552706 215076 552712
rect 214656 552016 214708 552022
rect 214656 551958 214708 551964
rect 214564 550248 214616 550254
rect 214564 550190 214616 550196
rect 215036 547963 215064 552706
rect 215772 547963 215800 552758
rect 215864 550202 215892 557506
rect 215956 550390 215984 630702
rect 216036 579692 216088 579698
rect 216036 579634 216088 579640
rect 216048 555694 216076 579634
rect 216680 564596 216732 564602
rect 216680 564538 216732 564544
rect 216692 557534 216720 564538
rect 216692 557506 217180 557534
rect 216036 555688 216088 555694
rect 216036 555630 216088 555636
rect 215944 550384 215996 550390
rect 215944 550326 215996 550332
rect 215864 550174 216444 550202
rect 216416 547963 216444 550174
rect 217152 547963 217180 557506
rect 217336 550458 217364 630974
rect 220176 630896 220228 630902
rect 220176 630838 220228 630844
rect 220084 630828 220136 630834
rect 220084 630770 220136 630776
rect 217416 627972 217468 627978
rect 217416 627914 217468 627920
rect 217428 554402 217456 627914
rect 218060 610020 218112 610026
rect 218060 609962 218112 609968
rect 217508 597576 217560 597582
rect 217508 597518 217560 597524
rect 217520 561202 217548 597518
rect 217508 561196 217560 561202
rect 217508 561138 217560 561144
rect 217416 554396 217468 554402
rect 217416 554338 217468 554344
rect 217876 552900 217928 552906
rect 217876 552842 217928 552848
rect 217324 550452 217376 550458
rect 217324 550394 217376 550400
rect 217888 547963 217916 552842
rect 218072 552786 218100 609962
rect 218152 572756 218204 572762
rect 218152 572698 218204 572704
rect 218164 557534 218192 572698
rect 219440 565276 219492 565282
rect 219440 565218 219492 565224
rect 218164 557506 219296 557534
rect 218072 552758 218652 552786
rect 218624 547963 218652 552758
rect 219268 547963 219296 557506
rect 219452 552838 219480 565218
rect 219440 552832 219492 552838
rect 219440 552774 219492 552780
rect 220096 550322 220124 630770
rect 220084 550316 220136 550322
rect 220084 550258 220136 550264
rect 219992 550248 220044 550254
rect 219992 550190 220044 550196
rect 220004 547963 220032 550190
rect 220188 550118 220216 630838
rect 220268 590708 220320 590714
rect 220268 590650 220320 590656
rect 220280 551682 220308 590650
rect 220360 569968 220412 569974
rect 220360 569910 220412 569916
rect 220372 564602 220400 569910
rect 220820 565140 220872 565146
rect 220820 565082 220872 565088
rect 220360 564596 220412 564602
rect 220360 564538 220412 564544
rect 220832 557534 220860 565082
rect 220832 557506 221504 557534
rect 220728 552832 220780 552838
rect 220728 552774 220780 552780
rect 220268 551676 220320 551682
rect 220268 551618 220320 551624
rect 220176 550112 220228 550118
rect 220176 550054 220228 550060
rect 220740 547963 220768 552774
rect 221476 547963 221504 557506
rect 222212 552838 222240 632878
rect 222844 615528 222896 615534
rect 222844 615470 222896 615476
rect 222292 565208 222344 565214
rect 222292 565150 222344 565156
rect 222200 552832 222252 552838
rect 222200 552774 222252 552780
rect 222304 548162 222332 565150
rect 222856 558482 222884 615470
rect 222844 558476 222896 558482
rect 222844 558418 222896 558424
rect 222844 552832 222896 552838
rect 222844 552774 222896 552780
rect 222228 548134 222332 548162
rect 222228 547944 222256 548134
rect 222856 547963 222884 552774
rect 223592 547963 223620 632946
rect 223672 612808 223724 612814
rect 223672 612750 223724 612756
rect 223684 557534 223712 612750
rect 223684 557506 224356 557534
rect 224328 547963 224356 557506
rect 226352 552786 226380 633966
rect 231124 633888 231176 633894
rect 231124 633830 231176 633836
rect 228364 631304 228416 631310
rect 228364 631246 228416 631252
rect 226432 576904 226484 576910
rect 226432 576846 226484 576852
rect 226444 557534 226472 576846
rect 227720 566704 227772 566710
rect 227720 566646 227772 566652
rect 226444 557506 227208 557534
rect 226352 552758 226472 552786
rect 225052 550316 225104 550322
rect 225052 550258 225104 550264
rect 225064 547963 225092 550258
rect 225788 550112 225840 550118
rect 225788 550054 225840 550060
rect 225800 547963 225828 550054
rect 226444 547963 226472 552758
rect 227180 547963 227208 557506
rect 227732 552838 227760 566646
rect 227812 565412 227864 565418
rect 227812 565354 227864 565360
rect 227824 557534 227852 565354
rect 227824 557506 227944 557534
rect 227720 552832 227772 552838
rect 227720 552774 227772 552780
rect 227916 547963 227944 557506
rect 228376 550186 228404 631246
rect 229744 600364 229796 600370
rect 229744 600306 229796 600312
rect 229284 554124 229336 554130
rect 229284 554066 229336 554072
rect 228640 552832 228692 552838
rect 228640 552774 228692 552780
rect 228364 550180 228416 550186
rect 228364 550122 228416 550128
rect 228652 547963 228680 552774
rect 229296 547963 229324 554066
rect 229756 551614 229784 600306
rect 230480 565480 230532 565486
rect 230480 565422 230532 565428
rect 230492 557534 230520 565422
rect 230492 557506 230980 557534
rect 229744 551608 229796 551614
rect 229744 551550 229796 551556
rect 230020 550588 230072 550594
rect 230020 550530 230072 550536
rect 230032 547963 230060 550530
rect 230756 550180 230808 550186
rect 230756 550122 230808 550128
rect 230768 547963 230796 550122
rect 230952 549930 230980 557506
rect 231136 550594 231164 633830
rect 234620 633820 234672 633826
rect 234620 633762 234672 633768
rect 233884 631236 233936 631242
rect 233884 631178 233936 631184
rect 231216 631100 231268 631106
rect 231216 631042 231268 631048
rect 231124 550588 231176 550594
rect 231124 550530 231176 550536
rect 231228 550050 231256 631042
rect 233240 622464 233292 622470
rect 233240 622406 233292 622412
rect 232504 619676 232556 619682
rect 232504 619618 232556 619624
rect 231860 587920 231912 587926
rect 231860 587862 231912 587868
rect 231872 552838 231900 587862
rect 231952 565344 232004 565350
rect 231952 565286 232004 565292
rect 231964 557534 231992 565286
rect 231964 557506 232268 557534
rect 231860 552832 231912 552838
rect 231860 552774 231912 552780
rect 231216 550044 231268 550050
rect 231216 549986 231268 549992
rect 230952 549902 231532 549930
rect 231504 547963 231532 549902
rect 232240 547963 232268 557506
rect 232516 557122 232544 619618
rect 233252 557534 233280 622406
rect 233252 557506 233648 557534
rect 232504 557116 232556 557122
rect 232504 557058 232556 557064
rect 232872 552832 232924 552838
rect 232872 552774 232924 552780
rect 232884 547963 232912 552774
rect 233620 547963 233648 557506
rect 233896 550254 233924 631178
rect 234632 557534 234660 633762
rect 235264 633616 235316 633622
rect 235264 633558 235316 633564
rect 234632 557506 235120 557534
rect 234344 550588 234396 550594
rect 234344 550530 234396 550536
rect 233884 550248 233936 550254
rect 233884 550190 233936 550196
rect 234356 547963 234384 550530
rect 235092 547963 235120 557506
rect 235276 553042 235304 633558
rect 235356 585200 235408 585206
rect 235356 585142 235408 585148
rect 235368 554198 235396 585142
rect 235448 565548 235500 565554
rect 235448 565490 235500 565496
rect 235356 554192 235408 554198
rect 235356 554134 235408 554140
rect 235264 553036 235316 553042
rect 235264 552978 235316 552984
rect 235460 550322 235488 565490
rect 236656 550594 236684 634170
rect 239404 634160 239456 634166
rect 239404 634102 239456 634108
rect 257068 634160 257120 634166
rect 257068 634102 257120 634108
rect 238208 634092 238260 634098
rect 238208 634034 238260 634040
rect 237380 633548 237432 633554
rect 237380 633490 237432 633496
rect 237392 629950 237420 633490
rect 237840 632732 237892 632738
rect 237840 632674 237892 632680
rect 237852 630698 237880 632674
rect 238116 631168 238168 631174
rect 238116 631110 238168 631116
rect 237840 630692 237892 630698
rect 237840 630634 237892 630640
rect 237380 629944 237432 629950
rect 237380 629886 237432 629892
rect 237378 628688 237434 628697
rect 237378 628623 237434 628632
rect 237392 627978 237420 628623
rect 237380 627972 237432 627978
rect 237380 627914 237432 627920
rect 237852 625154 237880 630634
rect 237852 625126 238064 625154
rect 237380 622464 237432 622470
rect 237378 622432 237380 622441
rect 237432 622432 237434 622441
rect 237378 622367 237434 622376
rect 237378 619712 237434 619721
rect 237378 619647 237380 619656
rect 237432 619647 237434 619656
rect 237380 619618 237432 619624
rect 237378 616312 237434 616321
rect 237378 616247 237434 616256
rect 237392 615534 237420 616247
rect 237380 615528 237432 615534
rect 237380 615470 237432 615476
rect 237378 613592 237434 613601
rect 237378 613527 237434 613536
rect 237392 612814 237420 613527
rect 237380 612808 237432 612814
rect 237380 612750 237432 612756
rect 237378 610192 237434 610201
rect 237378 610127 237434 610136
rect 237392 610026 237420 610127
rect 237380 610020 237432 610026
rect 237380 609962 237432 609968
rect 238036 604217 238064 625126
rect 238022 604208 238078 604217
rect 238022 604143 238078 604152
rect 237378 601352 237434 601361
rect 237378 601287 237434 601296
rect 237392 600370 237420 601287
rect 237380 600364 237432 600370
rect 237380 600306 237432 600312
rect 237378 597952 237434 597961
rect 237378 597887 237434 597896
rect 237392 597582 237420 597887
rect 237380 597576 237432 597582
rect 237380 597518 237432 597524
rect 237378 595232 237434 595241
rect 237378 595167 237434 595176
rect 237392 594862 237420 595167
rect 237380 594856 237432 594862
rect 237380 594798 237432 594804
rect 237378 591832 237434 591841
rect 237378 591767 237434 591776
rect 237392 590714 237420 591767
rect 237380 590708 237432 590714
rect 237380 590650 237432 590656
rect 237378 589112 237434 589121
rect 237378 589047 237434 589056
rect 237392 587926 237420 589047
rect 237380 587920 237432 587926
rect 237380 587862 237432 587868
rect 237378 585712 237434 585721
rect 237378 585647 237434 585656
rect 237392 585206 237420 585647
rect 237380 585200 237432 585206
rect 237380 585142 237432 585148
rect 236734 582992 236790 583001
rect 236734 582927 236790 582936
rect 236748 558414 236776 582927
rect 237378 579728 237434 579737
rect 237378 579663 237380 579672
rect 237432 579663 237434 579672
rect 237380 579634 237432 579640
rect 237380 576904 237432 576910
rect 237378 576872 237380 576881
rect 237432 576872 237434 576881
rect 237378 576807 237434 576816
rect 237378 573472 237434 573481
rect 237378 573407 237434 573416
rect 237392 572762 237420 573407
rect 237380 572756 237432 572762
rect 237380 572698 237432 572704
rect 237378 570752 237434 570761
rect 237378 570687 237434 570696
rect 237392 569974 237420 570687
rect 237380 569968 237432 569974
rect 237380 569910 237432 569916
rect 236736 558408 236788 558414
rect 236736 558350 236788 558356
rect 237932 552084 237984 552090
rect 237932 552026 237984 552032
rect 236644 550588 236696 550594
rect 236644 550530 236696 550536
rect 235448 550316 235500 550322
rect 235448 550258 235500 550264
rect 236460 548208 236512 548214
rect 236460 548150 236512 548156
rect 237194 548176 237250 548185
rect 235816 548140 235868 548146
rect 235816 548082 235868 548088
rect 235828 547963 235856 548082
rect 236472 547963 236500 548150
rect 237194 548111 237250 548120
rect 237208 547963 237236 548111
rect 237944 547963 237972 552026
rect 238128 549914 238156 631110
rect 238220 557054 238248 634034
rect 238944 632528 238996 632534
rect 238944 632470 238996 632476
rect 238852 627836 238904 627842
rect 238852 627778 238904 627784
rect 238298 625832 238354 625841
rect 238298 625767 238354 625776
rect 238208 557048 238260 557054
rect 238208 556990 238260 556996
rect 238312 551546 238340 625767
rect 238864 563922 238892 627778
rect 238956 607617 238984 632470
rect 239036 632324 239088 632330
rect 239036 632266 239088 632272
rect 238942 607608 238998 607617
rect 238942 607543 238998 607552
rect 238852 563916 238904 563922
rect 238852 563858 238904 563864
rect 239048 557534 239076 632266
rect 239416 561270 239444 634102
rect 251364 634092 251416 634098
rect 251364 634034 251416 634040
rect 248788 633888 248840 633894
rect 248788 633830 248840 633836
rect 239588 633752 239640 633758
rect 239588 633694 239640 633700
rect 239496 630692 239548 630698
rect 239496 630634 239548 630640
rect 239508 562630 239536 630634
rect 239600 563990 239628 633694
rect 245660 633684 245712 633690
rect 245660 633626 245712 633632
rect 245672 630986 245700 633626
rect 248800 630986 248828 633830
rect 249340 633684 249392 633690
rect 249340 633626 249392 633632
rect 249352 633010 249380 633626
rect 249340 633004 249392 633010
rect 249340 632946 249392 632952
rect 251376 630986 251404 634034
rect 254492 633548 254544 633554
rect 254492 633490 254544 633496
rect 254504 630986 254532 633490
rect 255320 633480 255372 633486
rect 255320 633422 255372 633428
rect 255332 632942 255360 633422
rect 255320 632936 255372 632942
rect 255320 632878 255372 632884
rect 257080 630986 257108 634102
rect 300308 634024 300360 634030
rect 300308 633966 300360 633972
rect 289268 633956 289320 633962
rect 289268 633898 289320 633904
rect 274640 633752 274692 633758
rect 274640 633694 274692 633700
rect 262956 633480 263008 633486
rect 262956 633422 263008 633428
rect 260380 631032 260432 631038
rect 245672 630958 245870 630986
rect 248800 630958 249090 630986
rect 251376 630958 251666 630986
rect 254504 630958 254886 630986
rect 257080 630958 257462 630986
rect 262968 630986 262996 633422
rect 266544 631236 266596 631242
rect 266544 631178 266596 631184
rect 260432 630980 260682 630986
rect 260380 630974 260682 630980
rect 260392 630958 260682 630974
rect 262968 630958 263258 630986
rect 266556 630850 266584 631178
rect 271972 631100 272024 631106
rect 271972 631042 272024 631048
rect 271984 630986 272012 631042
rect 274652 630986 274680 633694
rect 280252 631304 280304 631310
rect 280252 631246 280304 631252
rect 277676 631168 277728 631174
rect 277676 631110 277728 631116
rect 277688 630986 277716 631110
rect 280264 630986 280292 631246
rect 289280 630986 289308 633898
rect 295524 633684 295576 633690
rect 295524 633626 295576 633632
rect 291844 633616 291896 633622
rect 291844 633558 291896 633564
rect 291856 630986 291884 633558
rect 295536 630986 295564 633626
rect 268672 630970 269054 630986
rect 268660 630964 269054 630970
rect 268712 630958 269054 630964
rect 271984 630958 272274 630986
rect 274652 630958 274850 630986
rect 277688 630958 278070 630986
rect 280264 630958 280646 630986
rect 289280 630958 289662 630986
rect 291856 630958 292238 630986
rect 295458 630958 295564 630986
rect 300320 630986 300348 633966
rect 304264 633888 304316 633894
rect 304264 633830 304316 633836
rect 300320 630958 300610 630986
rect 268660 630906 268712 630912
rect 266478 630822 266584 630850
rect 283564 630896 283616 630902
rect 283616 630844 283866 630850
rect 283564 630838 283866 630844
rect 283576 630822 283866 630838
rect 286152 630834 286442 630850
rect 286140 630828 286442 630834
rect 286192 630822 286442 630828
rect 286140 630770 286192 630776
rect 297732 630760 297784 630766
rect 242912 630698 243294 630714
rect 297784 630708 298034 630714
rect 297732 630702 298034 630708
rect 242900 630692 243294 630698
rect 242952 630686 243294 630692
rect 297744 630686 298034 630702
rect 242900 630634 242952 630640
rect 239784 630414 240074 630442
rect 239784 627842 239812 630414
rect 300858 628144 300914 628153
rect 300858 628079 300914 628088
rect 239772 627836 239824 627842
rect 239772 627778 239824 627784
rect 288532 568404 288584 568410
rect 288532 568346 288584 568352
rect 287060 568268 287112 568274
rect 287060 568210 287112 568216
rect 266360 568200 266412 568206
rect 239784 568126 240074 568154
rect 241532 568126 242650 568154
rect 244292 568126 245226 568154
rect 248446 568126 248552 568154
rect 239784 565146 239812 568126
rect 239772 565140 239824 565146
rect 239772 565082 239824 565088
rect 239588 563984 239640 563990
rect 239588 563926 239640 563932
rect 239496 562624 239548 562630
rect 239496 562566 239548 562572
rect 239404 561264 239456 561270
rect 239404 561206 239456 561212
rect 240140 561128 240192 561134
rect 240140 561070 240192 561076
rect 240152 557534 240180 561070
rect 239048 557506 239444 557534
rect 240152 557506 240824 557534
rect 238300 551540 238352 551546
rect 238300 551482 238352 551488
rect 238116 549908 238168 549914
rect 238116 549850 238168 549856
rect 238666 549536 238722 549545
rect 238666 549471 238722 549480
rect 238680 547963 238708 549471
rect 239416 547963 239444 557506
rect 240048 548276 240100 548282
rect 240048 548218 240100 548224
rect 240060 547963 240088 548218
rect 240796 547963 240824 557506
rect 241532 550118 241560 568126
rect 242900 562556 242952 562562
rect 242900 562498 242952 562504
rect 241520 550112 241572 550118
rect 241520 550054 241572 550060
rect 242256 550112 242308 550118
rect 242256 550054 242308 550060
rect 241518 549672 241574 549681
rect 241518 549607 241574 549616
rect 241532 547963 241560 549607
rect 242268 547963 242296 550054
rect 242912 547963 242940 562498
rect 244292 559774 244320 568126
rect 248524 565554 248552 568126
rect 250640 568126 251022 568154
rect 253952 568126 254242 568154
rect 256818 568126 256924 568154
rect 248512 565548 248564 565554
rect 248512 565490 248564 565496
rect 249064 565548 249116 565554
rect 249064 565490 249116 565496
rect 244924 564460 244976 564466
rect 244924 564402 244976 564408
rect 244280 559768 244332 559774
rect 244280 559710 244332 559716
rect 244280 559632 244332 559638
rect 244280 559574 244332 559580
rect 244292 557534 244320 559574
rect 244292 557506 244596 557534
rect 244372 550656 244424 550662
rect 244372 550598 244424 550604
rect 243636 549500 243688 549506
rect 243636 549442 243688 549448
rect 243648 547963 243676 549442
rect 244384 547963 244412 550598
rect 244568 550066 244596 557506
rect 244936 550186 244964 564402
rect 246488 554192 246540 554198
rect 246488 554134 246540 554140
rect 244924 550180 244976 550186
rect 244924 550122 244976 550128
rect 244568 550038 245148 550066
rect 245120 547963 245148 550038
rect 245842 549944 245898 549953
rect 245842 549879 245898 549888
rect 245856 547963 245884 549879
rect 246500 547963 246528 554134
rect 247960 552832 248012 552838
rect 247960 552774 248012 552780
rect 247224 551336 247276 551342
rect 247224 551278 247276 551284
rect 247236 547963 247264 551278
rect 247972 547963 248000 552774
rect 249076 549982 249104 565490
rect 250640 564466 250668 568126
rect 250628 564460 250680 564466
rect 250628 564402 250680 564408
rect 251180 561196 251232 561202
rect 251180 561138 251232 561144
rect 249800 558408 249852 558414
rect 249800 558350 249852 558356
rect 249812 557534 249840 558350
rect 251192 557534 251220 561138
rect 252560 558272 252612 558278
rect 252560 558214 252612 558220
rect 252572 557534 252600 558214
rect 249812 557506 250116 557534
rect 251192 557506 251588 557534
rect 252572 557506 253704 557534
rect 249432 551472 249484 551478
rect 249432 551414 249484 551420
rect 249064 549976 249116 549982
rect 249064 549918 249116 549924
rect 248694 549808 248750 549817
rect 248694 549743 248750 549752
rect 248708 547963 248736 549743
rect 249444 547963 249472 551414
rect 250088 547963 250116 557506
rect 250812 556980 250864 556986
rect 250812 556922 250864 556928
rect 250824 547963 250852 556922
rect 251560 547963 251588 557506
rect 252928 552152 252980 552158
rect 252928 552094 252980 552100
rect 252284 549976 252336 549982
rect 252284 549918 252336 549924
rect 252296 547963 252324 549918
rect 252940 547963 252968 552094
rect 253676 547963 253704 557506
rect 253952 551410 253980 568126
rect 256896 567194 256924 568126
rect 259656 568126 260038 568154
rect 260840 568132 260892 568138
rect 258080 568064 258132 568070
rect 258080 568006 258132 568012
rect 256712 567166 256924 567194
rect 255320 562624 255372 562630
rect 255320 562566 255372 562572
rect 255332 552634 255360 562566
rect 256712 559842 256740 567166
rect 256700 559836 256752 559842
rect 256700 559778 256752 559784
rect 258092 557534 258120 568006
rect 259656 565486 259684 568126
rect 260840 568074 260892 568080
rect 262232 568126 262614 568154
rect 265544 568126 265834 568154
rect 266360 568142 266412 568148
rect 259644 565480 259696 565486
rect 259644 565422 259696 565428
rect 259460 565140 259512 565146
rect 259460 565082 259512 565088
rect 258092 557506 258764 557534
rect 257988 554260 258040 554266
rect 257988 554202 258040 554208
rect 255320 552628 255372 552634
rect 255320 552570 255372 552576
rect 256516 552628 256568 552634
rect 256516 552570 256568 552576
rect 253940 551404 253992 551410
rect 253940 551346 253992 551352
rect 255872 551200 255924 551206
rect 255872 551142 255924 551148
rect 255134 549400 255190 549409
rect 255134 549335 255190 549344
rect 254400 548140 254452 548146
rect 254400 548082 254452 548088
rect 254412 547963 254440 548082
rect 255148 547963 255176 549335
rect 255884 547963 255912 551142
rect 256528 547963 256556 552570
rect 257252 550248 257304 550254
rect 257252 550190 257304 550196
rect 257264 547963 257292 550190
rect 258000 547963 258028 554202
rect 258736 547963 258764 557506
rect 259472 547963 259500 565082
rect 260852 557534 260880 568074
rect 260852 557506 261616 557534
rect 260104 552968 260156 552974
rect 260104 552910 260156 552916
rect 260116 547963 260144 552910
rect 260840 548344 260892 548350
rect 260840 548286 260892 548292
rect 260852 547963 260880 548286
rect 261588 547963 261616 557506
rect 262232 554334 262260 568126
rect 265544 565418 265572 568126
rect 265532 565412 265584 565418
rect 265532 565354 265584 565360
rect 263600 563916 263652 563922
rect 263600 563858 263652 563864
rect 263612 557534 263640 563858
rect 263612 557506 263732 557534
rect 262220 554328 262272 554334
rect 262220 554270 262272 554276
rect 263048 550724 263100 550730
rect 263048 550666 263100 550672
rect 262312 548412 262364 548418
rect 262312 548354 262364 548360
rect 262324 547963 262352 548354
rect 263060 547963 263088 550666
rect 263704 547963 263732 557506
rect 266372 552634 266400 568142
rect 268120 568126 268410 568154
rect 271248 568126 271630 568154
rect 273824 568126 274206 568154
rect 277426 568126 277532 568154
rect 268120 565282 268148 568126
rect 269120 566772 269172 566778
rect 269120 566714 269172 566720
rect 268108 565276 268160 565282
rect 268108 565218 268160 565224
rect 266452 561264 266504 561270
rect 266452 561206 266504 561212
rect 266464 557534 266492 561206
rect 267740 558952 267792 558958
rect 267740 558894 267792 558900
rect 267752 557534 267780 558894
rect 266464 557506 266584 557534
rect 267752 557506 268056 557534
rect 266360 552628 266412 552634
rect 266360 552570 266412 552576
rect 265900 551268 265952 551274
rect 265900 551210 265952 551216
rect 265164 550996 265216 551002
rect 265164 550938 265216 550944
rect 264428 550792 264480 550798
rect 264428 550734 264480 550740
rect 264440 547963 264468 550734
rect 265176 547963 265204 550938
rect 265912 547963 265940 551210
rect 266556 547963 266584 557506
rect 267280 552628 267332 552634
rect 267280 552570 267332 552576
rect 267292 547963 267320 552570
rect 268028 547963 268056 557506
rect 269132 552786 269160 566714
rect 271248 565554 271276 568126
rect 271236 565548 271288 565554
rect 271236 565490 271288 565496
rect 269764 565480 269816 565486
rect 269764 565422 269816 565428
rect 269212 565276 269264 565282
rect 269212 565218 269264 565224
rect 269224 557534 269252 565218
rect 269224 557506 269620 557534
rect 269592 552786 269620 557506
rect 269776 552906 269804 565422
rect 273352 565412 273404 565418
rect 273352 565354 273404 565360
rect 273260 562692 273312 562698
rect 273260 562634 273312 562640
rect 270500 558476 270552 558482
rect 270500 558418 270552 558424
rect 270512 557534 270540 558418
rect 270512 557506 271644 557534
rect 269764 552900 269816 552906
rect 269764 552842 269816 552848
rect 269132 552758 269528 552786
rect 269592 552758 270172 552786
rect 268752 548616 268804 548622
rect 268752 548558 268804 548564
rect 268764 547963 268792 548558
rect 269500 547963 269528 552758
rect 270144 547963 270172 552758
rect 270868 550180 270920 550186
rect 270868 550122 270920 550128
rect 270880 547963 270908 550122
rect 271616 547963 271644 557506
rect 273272 552634 273300 562634
rect 273364 562494 273392 565354
rect 273824 565214 273852 568126
rect 273812 565208 273864 565214
rect 273812 565150 273864 565156
rect 273352 562488 273404 562494
rect 273352 562430 273404 562436
rect 277504 559706 277532 568126
rect 279712 568126 280002 568154
rect 282932 568126 283222 568154
rect 285798 568126 285904 568154
rect 279712 565350 279740 568126
rect 282932 565486 282960 568126
rect 285876 567194 285904 568126
rect 285692 567166 285904 567194
rect 282920 565480 282972 565486
rect 282920 565422 282972 565428
rect 279700 565344 279752 565350
rect 279700 565286 279752 565292
rect 280160 565208 280212 565214
rect 280160 565150 280212 565156
rect 277492 559700 277544 559706
rect 277492 559642 277544 559648
rect 280172 557534 280200 565150
rect 282184 564460 282236 564466
rect 282184 564402 282236 564408
rect 280172 557506 280936 557534
rect 279516 554328 279568 554334
rect 279516 554270 279568 554276
rect 275192 552900 275244 552906
rect 275192 552842 275244 552848
rect 273260 552628 273312 552634
rect 273260 552570 273312 552576
rect 274456 552628 274508 552634
rect 274456 552570 274508 552576
rect 273076 551132 273128 551138
rect 273076 551074 273128 551080
rect 272340 548480 272392 548486
rect 272340 548422 272392 548428
rect 272352 547963 272380 548422
rect 273088 547963 273116 551074
rect 273720 551064 273772 551070
rect 273720 551006 273772 551012
rect 273732 547963 273760 551006
rect 274468 547963 274496 552570
rect 275204 547963 275232 552842
rect 276572 549840 276624 549846
rect 276572 549782 276624 549788
rect 275928 549704 275980 549710
rect 275928 549646 275980 549652
rect 275940 547963 275968 549646
rect 276584 547963 276612 549782
rect 277308 549772 277360 549778
rect 277308 549714 277360 549720
rect 277320 547963 277348 549714
rect 278044 549296 278096 549302
rect 278044 549238 278096 549244
rect 278056 547963 278084 549238
rect 278780 548752 278832 548758
rect 278780 548694 278832 548700
rect 278792 547963 278820 548694
rect 279528 547963 279556 554270
rect 280160 549908 280212 549914
rect 280160 549850 280212 549856
rect 280172 547963 280200 549850
rect 280908 547963 280936 557506
rect 282196 555558 282224 564402
rect 285692 558346 285720 567166
rect 285680 558340 285732 558346
rect 285680 558282 285732 558288
rect 287072 557534 287100 568210
rect 287072 557506 288112 557534
rect 282368 555620 282420 555626
rect 282368 555562 282420 555568
rect 282184 555552 282236 555558
rect 282184 555494 282236 555500
rect 281632 548684 281684 548690
rect 281632 548626 281684 548632
rect 281644 547963 281672 548626
rect 282380 547963 282408 555562
rect 283748 555552 283800 555558
rect 283748 555494 283800 555500
rect 283104 549432 283156 549438
rect 283104 549374 283156 549380
rect 283116 547963 283144 549374
rect 283760 547963 283788 555494
rect 286692 552356 286744 552362
rect 286692 552298 286744 552304
rect 285220 552288 285272 552294
rect 285220 552230 285272 552236
rect 284484 549636 284536 549642
rect 284484 549578 284536 549584
rect 284496 547963 284524 549578
rect 285232 547963 285260 552230
rect 285956 552220 286008 552226
rect 285956 552162 286008 552168
rect 285968 547963 285996 552162
rect 286704 547963 286732 552298
rect 287336 550860 287388 550866
rect 287336 550802 287388 550808
rect 287348 547963 287376 550802
rect 287612 549500 287664 549506
rect 287612 549442 287664 549448
rect 287624 548554 287652 549442
rect 287888 549364 287940 549370
rect 287888 549306 287940 549312
rect 287900 548690 287928 549306
rect 287888 548684 287940 548690
rect 287888 548626 287940 548632
rect 287612 548548 287664 548554
rect 287612 548490 287664 548496
rect 288084 547963 288112 557506
rect 288544 553394 288572 568346
rect 288624 568336 288676 568342
rect 288624 568278 288676 568284
rect 288636 557534 288664 568278
rect 288728 568126 289018 568154
rect 291304 568126 291594 568154
rect 294432 568126 294814 568154
rect 297008 568126 297390 568154
rect 300320 568126 300610 568154
rect 288728 564466 288756 568126
rect 289820 567724 289872 567730
rect 289820 567666 289872 567672
rect 288716 564460 288768 564466
rect 288716 564402 288768 564408
rect 289832 557534 289860 567666
rect 291200 567656 291252 567662
rect 291200 567598 291252 567604
rect 288636 557506 289584 557534
rect 289832 557506 290228 557534
rect 288544 553366 288848 553394
rect 288820 547963 288848 553366
rect 289556 547963 289584 557506
rect 290200 547963 290228 557506
rect 290924 552424 290976 552430
rect 290924 552366 290976 552372
rect 290936 547963 290964 552366
rect 291212 550594 291240 567598
rect 291304 556850 291332 568126
rect 293960 567792 294012 567798
rect 293960 567734 294012 567740
rect 291844 565344 291896 565350
rect 291844 565286 291896 565292
rect 291292 556844 291344 556850
rect 291292 556786 291344 556792
rect 291856 554062 291884 565286
rect 291844 554056 291896 554062
rect 291844 553998 291896 554004
rect 293972 552634 294000 567734
rect 294432 562426 294460 568126
rect 297008 565418 297036 568126
rect 296996 565412 297048 565418
rect 296996 565354 297048 565360
rect 300320 565350 300348 568126
rect 300872 567866 300900 628079
rect 300950 625424 301006 625433
rect 300950 625359 301006 625368
rect 300860 567860 300912 567866
rect 300860 567802 300912 567808
rect 300964 566710 300992 625359
rect 302882 621208 302938 621217
rect 302882 621143 302938 621152
rect 301134 618488 301190 618497
rect 301134 618423 301190 618432
rect 301042 615632 301098 615641
rect 301042 615567 301098 615576
rect 300952 566704 301004 566710
rect 300952 566646 301004 566652
rect 300308 565344 300360 565350
rect 300308 565286 300360 565292
rect 294420 562420 294472 562426
rect 294420 562362 294472 562368
rect 301056 561066 301084 615567
rect 301148 567934 301176 618423
rect 301226 612776 301282 612785
rect 301226 612711 301282 612720
rect 301136 567928 301188 567934
rect 301136 567870 301188 567876
rect 301240 563786 301268 612711
rect 302422 608968 302478 608977
rect 302422 608903 302478 608912
rect 301318 600400 301374 600409
rect 301318 600335 301374 600344
rect 301228 563780 301280 563786
rect 301228 563722 301280 563728
rect 301044 561060 301096 561066
rect 301044 561002 301096 561008
rect 301332 552702 301360 600335
rect 301410 594008 301466 594017
rect 301410 593943 301466 593952
rect 301424 566574 301452 593943
rect 302238 588024 302294 588033
rect 302238 587959 302294 587968
rect 301502 581768 301558 581777
rect 301502 581703 301558 581712
rect 301412 566568 301464 566574
rect 301412 566510 301464 566516
rect 301516 563854 301544 581703
rect 301594 575648 301650 575657
rect 301594 575583 301650 575592
rect 301608 566506 301636 575583
rect 301686 570072 301742 570081
rect 301686 570007 301742 570016
rect 301596 566500 301648 566506
rect 301596 566442 301648 566448
rect 301504 563848 301556 563854
rect 301504 563790 301556 563796
rect 301700 560998 301728 570007
rect 302252 566642 302280 587959
rect 302330 578368 302386 578377
rect 302330 578303 302386 578312
rect 302344 568002 302372 578303
rect 302332 567996 302384 568002
rect 302332 567938 302384 567944
rect 302240 566636 302292 566642
rect 302240 566578 302292 566584
rect 301688 560992 301740 560998
rect 301688 560934 301740 560940
rect 302436 555490 302464 608903
rect 302514 603120 302570 603129
rect 302514 603055 302570 603064
rect 302424 555484 302476 555490
rect 302424 555426 302476 555432
rect 302528 552770 302556 603055
rect 302700 596828 302752 596834
rect 302700 596770 302752 596776
rect 302712 596737 302740 596770
rect 302698 596728 302754 596737
rect 302698 596663 302754 596672
rect 302606 590744 302662 590753
rect 302606 590679 302662 590688
rect 302620 559570 302648 590679
rect 302712 568478 302740 596663
rect 302790 584488 302846 584497
rect 302790 584423 302846 584432
rect 302700 568472 302752 568478
rect 302700 568414 302752 568420
rect 302608 559564 302660 559570
rect 302608 559506 302660 559512
rect 302516 552764 302568 552770
rect 302516 552706 302568 552712
rect 301320 552696 301372 552702
rect 301320 552638 301372 552644
rect 293960 552628 294012 552634
rect 293960 552570 294012 552576
rect 295248 552628 295300 552634
rect 295248 552570 295300 552576
rect 293132 552492 293184 552498
rect 293132 552434 293184 552440
rect 291660 550928 291712 550934
rect 291660 550870 291712 550876
rect 291200 550588 291252 550594
rect 291200 550530 291252 550536
rect 291672 547963 291700 550870
rect 292396 550588 292448 550594
rect 292396 550530 292448 550536
rect 292408 547963 292436 550530
rect 293144 547963 293172 552434
rect 293960 549976 294012 549982
rect 293960 549918 294012 549924
rect 293972 548690 294000 549918
rect 294512 549568 294564 549574
rect 294512 549510 294564 549516
rect 293960 548684 294012 548690
rect 293960 548626 294012 548632
rect 293774 548176 293830 548185
rect 293774 548111 293830 548120
rect 293788 547963 293816 548111
rect 294524 547963 294552 549510
rect 295260 547963 295288 552570
rect 301504 551472 301556 551478
rect 301504 551414 301556 551420
rect 299572 550588 299624 550594
rect 299572 550530 299624 550536
rect 298836 550520 298888 550526
rect 298836 550462 298888 550468
rect 298098 550216 298154 550225
rect 298098 550151 298154 550160
rect 297362 550080 297418 550089
rect 297362 550015 297418 550024
rect 295984 549500 296036 549506
rect 295984 549442 296036 549448
rect 295996 547963 296024 549442
rect 296720 548820 296772 548826
rect 296720 548762 296772 548768
rect 296732 547963 296760 548762
rect 297376 547963 297404 550015
rect 298112 547963 298140 550151
rect 298848 547963 298876 550462
rect 299584 547963 299612 550530
rect 300584 550248 300636 550254
rect 300584 550190 300636 550196
rect 300124 549840 300176 549846
rect 300124 549782 300176 549788
rect 300136 521218 300164 549782
rect 300400 549772 300452 549778
rect 300400 549714 300452 549720
rect 300308 549296 300360 549302
rect 300308 549238 300360 549244
rect 300216 548616 300268 548622
rect 300216 548558 300268 548564
rect 300124 521212 300176 521218
rect 300124 521154 300176 521160
rect 300228 520062 300256 548558
rect 300320 521354 300348 549238
rect 300412 522918 300440 549714
rect 300492 549364 300544 549370
rect 300492 549306 300544 549312
rect 300504 522986 300532 549306
rect 300492 522980 300544 522986
rect 300492 522922 300544 522928
rect 300400 522912 300452 522918
rect 300400 522854 300452 522860
rect 300596 522850 300624 550190
rect 300768 548752 300820 548758
rect 300768 548694 300820 548700
rect 300780 542366 300808 548694
rect 300768 542360 300820 542366
rect 300768 542302 300820 542308
rect 300584 522844 300636 522850
rect 300584 522786 300636 522792
rect 300308 521348 300360 521354
rect 300308 521290 300360 521296
rect 301516 520169 301544 551414
rect 301596 551336 301648 551342
rect 301596 551278 301648 551284
rect 301502 520160 301558 520169
rect 301502 520095 301558 520104
rect 300216 520056 300268 520062
rect 300216 519998 300268 520004
rect 301608 519790 301636 551278
rect 301688 549908 301740 549914
rect 301688 549850 301740 549856
rect 301700 521286 301728 549850
rect 301778 549808 301834 549817
rect 301778 549743 301834 549752
rect 301792 522782 301820 549743
rect 301962 549672 302018 549681
rect 301962 549607 302018 549616
rect 301870 547904 301926 547913
rect 301870 547839 301926 547848
rect 301780 522776 301832 522782
rect 301780 522718 301832 522724
rect 301884 522714 301912 547839
rect 301872 522708 301924 522714
rect 301872 522650 301924 522656
rect 301976 522481 302004 549607
rect 302056 548208 302108 548214
rect 302056 548150 302108 548156
rect 302068 536790 302096 548150
rect 302606 540424 302662 540433
rect 302606 540359 302662 540368
rect 302620 539646 302648 540359
rect 302608 539640 302660 539646
rect 302608 539582 302660 539588
rect 302056 536784 302108 536790
rect 302056 536726 302108 536732
rect 301962 522472 302018 522481
rect 301962 522407 302018 522416
rect 301688 521280 301740 521286
rect 301688 521222 301740 521228
rect 301596 519784 301648 519790
rect 301596 519726 301648 519732
rect 57886 517984 57942 517993
rect 57886 517919 57942 517928
rect 57900 517546 57928 517919
rect 52368 517540 52420 517546
rect 52368 517482 52420 517488
rect 57888 517540 57940 517546
rect 57888 517482 57940 517488
rect 51908 486532 51960 486538
rect 51908 486474 51960 486480
rect 51816 485240 51868 485246
rect 51816 485182 51868 485188
rect 45468 485172 45520 485178
rect 45468 485114 45520 485120
rect 43902 482352 43958 482361
rect 43902 482287 43958 482296
rect 42614 480040 42670 480049
rect 42614 479975 42670 479984
rect 42524 479868 42576 479874
rect 42524 479810 42576 479816
rect 42432 479800 42484 479806
rect 42432 479742 42484 479748
rect 42340 479664 42392 479670
rect 42340 479606 42392 479612
rect 42248 467288 42300 467294
rect 42248 467230 42300 467236
rect 41328 467220 41380 467226
rect 41328 467162 41380 467168
rect 41340 166326 41368 467162
rect 42156 465860 42208 465866
rect 42156 465802 42208 465808
rect 42168 377126 42196 465802
rect 42156 377120 42208 377126
rect 42156 377062 42208 377068
rect 42260 271794 42288 467230
rect 42352 273222 42380 479606
rect 42340 273216 42392 273222
rect 42340 273158 42392 273164
rect 42444 272882 42472 479742
rect 42432 272876 42484 272882
rect 42432 272818 42484 272824
rect 42248 271788 42300 271794
rect 42248 271730 42300 271736
rect 42536 271726 42564 479810
rect 42524 271720 42576 271726
rect 42524 271662 42576 271668
rect 41328 166320 41380 166326
rect 41328 166262 41380 166268
rect 21364 97980 21416 97986
rect 21364 97922 21416 97928
rect 42628 70378 42656 479975
rect 43718 477184 43774 477193
rect 43718 477119 43774 477128
rect 43534 476912 43590 476921
rect 43534 476847 43590 476856
rect 43444 472660 43496 472666
rect 43444 472602 43496 472608
rect 43352 468512 43404 468518
rect 43352 468454 43404 468460
rect 43260 465996 43312 466002
rect 43260 465938 43312 465944
rect 42708 465724 42760 465730
rect 42708 465666 42760 465672
rect 42616 70372 42668 70378
rect 42616 70314 42668 70320
rect 42720 56302 42748 465666
rect 43272 378146 43300 465938
rect 43260 378140 43312 378146
rect 43260 378082 43312 378088
rect 43364 273630 43392 468454
rect 43352 273624 43404 273630
rect 43352 273566 43404 273572
rect 43456 271862 43484 472602
rect 43444 271856 43496 271862
rect 43444 271798 43496 271804
rect 43548 268530 43576 476847
rect 43626 476776 43682 476785
rect 43626 476711 43682 476720
rect 43640 268666 43668 476711
rect 43628 268660 43680 268666
rect 43628 268602 43680 268608
rect 43536 268524 43588 268530
rect 43536 268466 43588 268472
rect 43732 268462 43760 477119
rect 43810 477048 43866 477057
rect 43810 476983 43866 476992
rect 43824 268598 43852 476983
rect 43812 268592 43864 268598
rect 43812 268534 43864 268540
rect 43720 268456 43772 268462
rect 43720 268398 43772 268404
rect 43916 267714 43944 482287
rect 43996 476944 44048 476950
rect 43996 476886 44048 476892
rect 44008 379098 44036 476886
rect 45008 476876 45060 476882
rect 45008 476818 45060 476824
rect 44732 476808 44784 476814
rect 44732 476750 44784 476756
rect 44088 467356 44140 467362
rect 44088 467298 44140 467304
rect 43996 379092 44048 379098
rect 43996 379034 44048 379040
rect 43994 378856 44050 378865
rect 43994 378791 44050 378800
rect 43904 267708 43956 267714
rect 43904 267650 43956 267656
rect 44008 57798 44036 378791
rect 43996 57792 44048 57798
rect 43996 57734 44048 57740
rect 44100 57526 44128 467298
rect 44640 416832 44692 416838
rect 44640 416774 44692 416780
rect 44652 375766 44680 416774
rect 44744 391950 44772 476750
rect 44916 471232 44968 471238
rect 44916 471174 44968 471180
rect 44824 471164 44876 471170
rect 44824 471106 44876 471112
rect 44732 391944 44784 391950
rect 44732 391886 44784 391892
rect 44836 378826 44864 471106
rect 44928 379030 44956 471174
rect 45020 380186 45048 476818
rect 45376 474564 45428 474570
rect 45376 474506 45428 474512
rect 45284 474088 45336 474094
rect 45284 474030 45336 474036
rect 45192 472796 45244 472802
rect 45192 472738 45244 472744
rect 45100 472728 45152 472734
rect 45100 472670 45152 472676
rect 45008 380180 45060 380186
rect 45008 380122 45060 380128
rect 44916 379024 44968 379030
rect 44916 378966 44968 378972
rect 44824 378820 44876 378826
rect 44824 378762 44876 378768
rect 44640 375760 44692 375766
rect 44640 375702 44692 375708
rect 45112 273562 45140 472670
rect 45100 273556 45152 273562
rect 45100 273498 45152 273504
rect 45204 273426 45232 472738
rect 45192 273420 45244 273426
rect 45192 273362 45244 273368
rect 45296 273290 45324 474030
rect 45388 273358 45416 474506
rect 45480 273494 45508 485114
rect 50436 482996 50488 483002
rect 50436 482938 50488 482944
rect 48044 482860 48096 482866
rect 48044 482802 48096 482808
rect 46664 482724 46716 482730
rect 46664 482666 46716 482672
rect 46570 482624 46626 482633
rect 46388 482588 46440 482594
rect 46570 482559 46626 482568
rect 46388 482530 46440 482536
rect 46296 482452 46348 482458
rect 46296 482394 46348 482400
rect 46112 479596 46164 479602
rect 46112 479538 46164 479544
rect 46020 464296 46072 464302
rect 46020 464238 46072 464244
rect 46032 418130 46060 464238
rect 46020 418124 46072 418130
rect 46020 418066 46072 418072
rect 46124 389094 46152 479538
rect 46204 477012 46256 477018
rect 46204 476954 46256 476960
rect 46112 389088 46164 389094
rect 46112 389030 46164 389036
rect 46216 379166 46244 476954
rect 46204 379160 46256 379166
rect 46204 379102 46256 379108
rect 46204 379024 46256 379030
rect 46204 378966 46256 378972
rect 46216 378214 46244 378966
rect 46204 378208 46256 378214
rect 46204 378150 46256 378156
rect 46216 287054 46244 378150
rect 46308 303618 46336 482394
rect 46296 303612 46348 303618
rect 46296 303554 46348 303560
rect 46400 300830 46428 482530
rect 46478 482488 46534 482497
rect 46478 482423 46534 482432
rect 46388 300824 46440 300830
rect 46388 300766 46440 300772
rect 46216 287026 46428 287054
rect 45468 273488 45520 273494
rect 45468 273430 45520 273436
rect 45376 273352 45428 273358
rect 45376 273294 45428 273300
rect 45284 273284 45336 273290
rect 45284 273226 45336 273232
rect 46020 273216 46072 273222
rect 46020 273158 46072 273164
rect 46032 272513 46060 273158
rect 46018 272504 46074 272513
rect 46018 272439 46074 272448
rect 46032 267734 46060 272439
rect 46400 271946 46428 287026
rect 46492 272202 46520 482423
rect 46480 272196 46532 272202
rect 46480 272138 46532 272144
rect 46584 272134 46612 482559
rect 46676 272406 46704 482666
rect 46756 482384 46808 482390
rect 46756 482326 46808 482332
rect 46664 272400 46716 272406
rect 46664 272342 46716 272348
rect 46572 272128 46624 272134
rect 46572 272070 46624 272076
rect 46400 271918 46612 271946
rect 46584 271017 46612 271918
rect 46570 271008 46626 271017
rect 46570 270943 46626 270952
rect 46480 268660 46532 268666
rect 46480 268602 46532 268608
rect 46388 268592 46440 268598
rect 46388 268534 46440 268540
rect 46204 268524 46256 268530
rect 46204 268466 46256 268472
rect 46032 267706 46152 267734
rect 46124 148578 46152 267706
rect 46216 165714 46244 268466
rect 46296 268456 46348 268462
rect 46296 268398 46348 268404
rect 46204 165708 46256 165714
rect 46204 165650 46256 165656
rect 46308 163606 46336 268398
rect 46296 163600 46348 163606
rect 46296 163542 46348 163548
rect 46400 162790 46428 268534
rect 46492 162858 46520 268602
rect 46480 162852 46532 162858
rect 46480 162794 46532 162800
rect 46388 162784 46440 162790
rect 46388 162726 46440 162732
rect 46584 148850 46612 270943
rect 46572 148844 46624 148850
rect 46572 148786 46624 148792
rect 46112 148572 46164 148578
rect 46112 148514 46164 148520
rect 46676 145382 46704 272342
rect 46768 271454 46796 482326
rect 47400 480140 47452 480146
rect 47400 480082 47452 480088
rect 46848 477420 46900 477426
rect 46848 477362 46900 477368
rect 46756 271448 46808 271454
rect 46756 271390 46808 271396
rect 46860 251190 46888 477362
rect 47412 269074 47440 480082
rect 47860 477148 47912 477154
rect 47860 477090 47912 477096
rect 47768 471096 47820 471102
rect 47768 471038 47820 471044
rect 47676 468444 47728 468450
rect 47676 468386 47728 468392
rect 47584 414044 47636 414050
rect 47584 413986 47636 413992
rect 47492 412684 47544 412690
rect 47492 412626 47544 412632
rect 47504 380866 47532 412626
rect 47492 380860 47544 380866
rect 47492 380802 47544 380808
rect 47596 380089 47624 413986
rect 47582 380080 47638 380089
rect 47582 380015 47638 380024
rect 47688 379273 47716 468386
rect 47780 379409 47808 471038
rect 47766 379400 47822 379409
rect 47766 379335 47822 379344
rect 47674 379264 47730 379273
rect 47674 379199 47730 379208
rect 47582 378992 47638 379001
rect 47582 378927 47638 378936
rect 47596 287054 47624 378927
rect 47688 373994 47716 379199
rect 47780 379001 47808 379335
rect 47766 378992 47822 379001
rect 47766 378927 47822 378936
rect 47872 378758 47900 477090
rect 47952 467152 48004 467158
rect 47952 467094 48004 467100
rect 47860 378752 47912 378758
rect 47860 378694 47912 378700
rect 47688 373966 47808 373994
rect 47780 287054 47808 373966
rect 47596 287026 47716 287054
rect 47780 287026 47900 287054
rect 47688 271561 47716 287026
rect 47674 271552 47730 271561
rect 47674 271487 47730 271496
rect 47400 269068 47452 269074
rect 47400 269010 47452 269016
rect 47584 268388 47636 268394
rect 47584 268330 47636 268336
rect 47596 267714 47624 268330
rect 47688 267734 47716 271487
rect 47872 271425 47900 287026
rect 47858 271416 47914 271425
rect 47858 271351 47914 271360
rect 47872 270314 47900 271351
rect 47964 270502 47992 467094
rect 48056 272610 48084 482802
rect 48136 482792 48188 482798
rect 48136 482734 48188 482740
rect 48148 272814 48176 482734
rect 49056 482520 49108 482526
rect 49056 482462 49108 482468
rect 48964 480004 49016 480010
rect 48964 479946 49016 479952
rect 48872 479732 48924 479738
rect 48872 479674 48924 479680
rect 48780 477080 48832 477086
rect 48780 477022 48832 477028
rect 48228 411324 48280 411330
rect 48228 411266 48280 411272
rect 48240 380798 48268 411266
rect 48228 380792 48280 380798
rect 48228 380734 48280 380740
rect 48792 380390 48820 477022
rect 48780 380384 48832 380390
rect 48780 380326 48832 380332
rect 48884 379370 48912 479674
rect 48872 379364 48924 379370
rect 48872 379306 48924 379312
rect 48872 378820 48924 378826
rect 48872 378762 48924 378768
rect 48884 378282 48912 378762
rect 48872 378276 48924 378282
rect 48872 378218 48924 378224
rect 48136 272808 48188 272814
rect 48136 272750 48188 272756
rect 48044 272604 48096 272610
rect 48044 272546 48096 272552
rect 47952 270496 48004 270502
rect 47952 270438 48004 270444
rect 47872 270286 48084 270314
rect 47584 267708 47636 267714
rect 47688 267706 47900 267734
rect 47584 267650 47636 267656
rect 46848 251184 46900 251190
rect 46848 251126 46900 251132
rect 46664 145376 46716 145382
rect 46664 145318 46716 145324
rect 47596 144702 47624 267650
rect 47872 148782 47900 267706
rect 47860 148776 47912 148782
rect 47860 148718 47912 148724
rect 48056 146266 48084 270286
rect 48044 146260 48096 146266
rect 48044 146202 48096 146208
rect 48148 145450 48176 272750
rect 48884 272218 48912 378218
rect 48976 272678 49004 479946
rect 48964 272672 49016 272678
rect 48964 272614 49016 272620
rect 49068 272474 49096 482462
rect 49148 479936 49200 479942
rect 49148 479878 49200 479884
rect 49056 272468 49108 272474
rect 49056 272410 49108 272416
rect 48884 272190 49096 272218
rect 48964 272128 49016 272134
rect 48964 272070 49016 272076
rect 48976 271998 49004 272070
rect 48964 271992 49016 271998
rect 48964 271934 49016 271940
rect 48228 271924 48280 271930
rect 48228 271866 48280 271872
rect 48240 147626 48268 271866
rect 48976 163742 49004 271934
rect 49068 271697 49096 272190
rect 49054 271688 49110 271697
rect 49054 271623 49110 271632
rect 48964 163736 49016 163742
rect 48964 163678 49016 163684
rect 49068 148714 49096 271623
rect 49160 251122 49188 479878
rect 50160 477216 50212 477222
rect 50160 477158 50212 477164
rect 49424 471572 49476 471578
rect 49424 471514 49476 471520
rect 49332 468648 49384 468654
rect 49332 468590 49384 468596
rect 49240 468580 49292 468586
rect 49240 468522 49292 468528
rect 49148 251116 49200 251122
rect 49148 251058 49200 251064
rect 49252 165481 49280 468522
rect 49238 165472 49294 165481
rect 49238 165407 49294 165416
rect 49344 165345 49372 468590
rect 49436 166938 49464 471514
rect 49514 471200 49570 471209
rect 49514 471135 49570 471144
rect 49424 166932 49476 166938
rect 49424 166874 49476 166880
rect 49330 165336 49386 165345
rect 49330 165271 49386 165280
rect 49528 165209 49556 471135
rect 49608 469124 49660 469130
rect 49608 469066 49660 469072
rect 49514 165200 49570 165209
rect 49514 165135 49570 165144
rect 49056 148708 49108 148714
rect 49056 148650 49108 148656
rect 48228 147620 48280 147626
rect 48228 147562 48280 147568
rect 48136 145444 48188 145450
rect 48136 145386 48188 145392
rect 47584 144696 47636 144702
rect 47584 144638 47636 144644
rect 49620 58818 49648 469066
rect 50172 379030 50200 477158
rect 50344 474292 50396 474298
rect 50344 474234 50396 474240
rect 50252 409896 50304 409902
rect 50252 409838 50304 409844
rect 50264 380662 50292 409838
rect 50252 380656 50304 380662
rect 50252 380598 50304 380604
rect 50160 379024 50212 379030
rect 50160 378966 50212 378972
rect 50158 273048 50214 273057
rect 50158 272983 50214 272992
rect 50068 272468 50120 272474
rect 50068 272410 50120 272416
rect 50080 272338 50108 272410
rect 50068 272332 50120 272338
rect 50068 272274 50120 272280
rect 50080 145654 50108 272274
rect 50172 163810 50200 272983
rect 50250 272912 50306 272921
rect 50250 272847 50306 272856
rect 50264 272678 50292 272847
rect 50252 272672 50304 272678
rect 50252 272614 50304 272620
rect 50160 163804 50212 163810
rect 50160 163746 50212 163752
rect 50068 145648 50120 145654
rect 50264 145625 50292 272614
rect 50356 271046 50384 474234
rect 50448 272746 50476 482938
rect 50528 482928 50580 482934
rect 50528 482870 50580 482876
rect 50436 272740 50488 272746
rect 50436 272682 50488 272688
rect 50540 272542 50568 482870
rect 50620 482656 50672 482662
rect 50620 482598 50672 482604
rect 50528 272536 50580 272542
rect 50528 272478 50580 272484
rect 50344 271040 50396 271046
rect 50344 270982 50396 270988
rect 50632 269754 50660 482598
rect 51632 482248 51684 482254
rect 51632 482190 51684 482196
rect 51540 474224 51592 474230
rect 51540 474166 51592 474172
rect 50896 471980 50948 471986
rect 50896 471922 50948 471928
rect 50804 471844 50856 471850
rect 50804 471786 50856 471792
rect 50712 471640 50764 471646
rect 50712 471582 50764 471588
rect 50620 269748 50672 269754
rect 50620 269690 50672 269696
rect 50724 166870 50752 471582
rect 50816 167006 50844 471786
rect 50804 167000 50856 167006
rect 50804 166942 50856 166948
rect 50712 166864 50764 166870
rect 50712 166806 50764 166812
rect 50908 164762 50936 471922
rect 51448 471776 51500 471782
rect 51448 471718 51500 471724
rect 51356 469192 51408 469198
rect 51356 469134 51408 469140
rect 51368 465050 51396 469134
rect 51460 465798 51488 471718
rect 51448 465792 51500 465798
rect 51448 465734 51500 465740
rect 51356 465044 51408 465050
rect 51356 464986 51408 464992
rect 50988 408536 51040 408542
rect 50988 408478 51040 408484
rect 51000 380769 51028 408478
rect 50986 380760 51042 380769
rect 50986 380695 51042 380704
rect 50986 379536 51042 379545
rect 50986 379471 51042 379480
rect 50896 164756 50948 164762
rect 50896 164698 50948 164704
rect 50896 162852 50948 162858
rect 50896 162794 50948 162800
rect 50908 162178 50936 162794
rect 50896 162172 50948 162178
rect 50896 162114 50948 162120
rect 50068 145590 50120 145596
rect 50250 145616 50306 145625
rect 50250 145551 50306 145560
rect 49608 58812 49660 58818
rect 49608 58754 49660 58760
rect 44088 57520 44140 57526
rect 44088 57462 44140 57468
rect 42708 56296 42760 56302
rect 42708 56238 42760 56244
rect 50908 55214 50936 162114
rect 51000 58750 51028 379471
rect 51448 272196 51500 272202
rect 51448 272138 51500 272144
rect 51460 163878 51488 272138
rect 51552 271318 51580 474166
rect 51644 272678 51672 482190
rect 51724 480208 51776 480214
rect 51724 480150 51776 480156
rect 51632 272672 51684 272678
rect 51632 272614 51684 272620
rect 51630 271824 51686 271833
rect 51630 271759 51686 271768
rect 51540 271312 51592 271318
rect 51540 271254 51592 271260
rect 51448 163872 51500 163878
rect 51448 163814 51500 163820
rect 50988 58744 51040 58750
rect 50988 58686 51040 58692
rect 51644 57866 51672 271759
rect 51736 270366 51764 480150
rect 51828 271182 51856 485182
rect 51816 271176 51868 271182
rect 51816 271118 51868 271124
rect 51920 271114 51948 486474
rect 52092 468784 52144 468790
rect 52092 468726 52144 468732
rect 52000 466404 52052 466410
rect 52000 466346 52052 466352
rect 52012 465225 52040 466346
rect 51998 465216 52054 465225
rect 51998 465151 52054 465160
rect 52000 465044 52052 465050
rect 52000 464986 52052 464992
rect 51908 271108 51960 271114
rect 51908 271050 51960 271056
rect 51724 270360 51776 270366
rect 51724 270302 51776 270308
rect 51736 267734 51764 270302
rect 51736 267706 51856 267734
rect 51724 146260 51776 146266
rect 51724 146202 51776 146208
rect 51736 145518 51764 146202
rect 51724 145512 51776 145518
rect 51724 145454 51776 145460
rect 51632 57860 51684 57866
rect 51632 57802 51684 57808
rect 51736 57254 51764 145454
rect 51828 144838 51856 267706
rect 52012 164898 52040 464986
rect 52104 165034 52132 468726
rect 52276 465928 52328 465934
rect 52276 465870 52328 465876
rect 52184 465792 52236 465798
rect 52184 465734 52236 465740
rect 52196 166734 52224 465734
rect 52184 166728 52236 166734
rect 52184 166670 52236 166676
rect 52184 165708 52236 165714
rect 52184 165650 52236 165656
rect 52092 165028 52144 165034
rect 52092 164970 52144 164976
rect 52000 164892 52052 164898
rect 52000 164834 52052 164840
rect 52092 162784 52144 162790
rect 52092 162726 52144 162732
rect 52104 162246 52132 162726
rect 52092 162240 52144 162246
rect 52092 162182 52144 162188
rect 52000 148708 52052 148714
rect 52000 148650 52052 148656
rect 51816 144832 51868 144838
rect 51816 144774 51868 144780
rect 51724 57248 51776 57254
rect 51724 57190 51776 57196
rect 52012 56030 52040 148650
rect 52104 56438 52132 162182
rect 52092 56432 52144 56438
rect 52092 56374 52144 56380
rect 52000 56024 52052 56030
rect 52000 55966 52052 55972
rect 50896 55208 50948 55214
rect 50896 55150 50948 55156
rect 52196 55078 52224 165650
rect 52288 59430 52316 465870
rect 52380 389162 52408 517482
rect 302712 510513 302740 568414
rect 302804 562358 302832 584423
rect 302792 562352 302844 562358
rect 302792 562294 302844 562300
rect 302896 556918 302924 621143
rect 302974 606384 303030 606393
rect 302974 606319 303030 606328
rect 302988 558210 303016 606319
rect 303066 572792 303122 572801
rect 303066 572727 303122 572736
rect 302976 558204 303028 558210
rect 302976 558146 303028 558152
rect 302884 556912 302936 556918
rect 302884 556854 302936 556860
rect 303080 554130 303108 572727
rect 303068 554124 303120 554130
rect 303068 554066 303120 554072
rect 304276 550526 304304 633830
rect 304356 633752 304408 633758
rect 304356 633694 304408 633700
rect 304368 550594 304396 633694
rect 304448 551200 304500 551206
rect 304448 551142 304500 551148
rect 304356 550588 304408 550594
rect 304356 550530 304408 550536
rect 304264 550520 304316 550526
rect 304264 550462 304316 550468
rect 302884 549704 302936 549710
rect 302884 549646 302936 549652
rect 302896 520810 302924 549646
rect 304264 548480 304316 548486
rect 304264 548422 304316 548428
rect 302976 548276 303028 548282
rect 302976 548218 303028 548224
rect 302988 527134 303016 548218
rect 302976 527128 303028 527134
rect 302976 527070 303028 527076
rect 302974 525464 303030 525473
rect 302974 525399 303030 525408
rect 302884 520804 302936 520810
rect 302884 520746 302936 520752
rect 302988 518226 303016 525399
rect 304276 519518 304304 548422
rect 304264 519512 304316 519518
rect 304264 519454 304316 519460
rect 304460 519450 304488 551142
rect 305656 520878 305684 700402
rect 364352 638246 364380 702406
rect 429856 700466 429884 703520
rect 429844 700460 429896 700466
rect 429844 700402 429896 700408
rect 434720 700460 434772 700466
rect 434720 700402 434772 700408
rect 405740 641028 405792 641034
rect 405740 640970 405792 640976
rect 318156 638240 318208 638246
rect 318156 638182 318208 638188
rect 364340 638240 364392 638246
rect 364340 638182 364392 638188
rect 307024 635792 307076 635798
rect 307024 635734 307076 635740
rect 305736 589348 305788 589354
rect 305736 589290 305788 589296
rect 305748 555626 305776 589290
rect 307036 561270 307064 635734
rect 318064 635588 318116 635594
rect 318064 635530 318116 635536
rect 316776 635384 316828 635390
rect 316776 635326 316828 635332
rect 313924 635180 313976 635186
rect 313924 635122 313976 635128
rect 309784 626612 309836 626618
rect 309784 626554 309836 626560
rect 307116 603152 307168 603158
rect 307116 603094 307168 603100
rect 307024 561264 307076 561270
rect 307024 561206 307076 561212
rect 307128 558414 307156 603094
rect 307208 597576 307260 597582
rect 307208 597518 307260 597524
rect 307220 565282 307248 597518
rect 307300 583772 307352 583778
rect 307300 583714 307352 583720
rect 307312 568546 307340 583714
rect 307300 568540 307352 568546
rect 307300 568482 307352 568488
rect 307208 565276 307260 565282
rect 307208 565218 307260 565224
rect 309796 558482 309824 626554
rect 311164 622464 311216 622470
rect 311164 622406 311216 622412
rect 309784 558476 309836 558482
rect 309784 558418 309836 558424
rect 307116 558408 307168 558414
rect 307116 558350 307168 558356
rect 305736 555620 305788 555626
rect 305736 555562 305788 555568
rect 311176 554334 311204 622406
rect 312544 612808 312596 612814
rect 312544 612750 312596 612756
rect 311256 574116 311308 574122
rect 311256 574058 311308 574064
rect 311164 554328 311216 554334
rect 311164 554270 311216 554276
rect 311268 552974 311296 574058
rect 312556 554198 312584 612750
rect 312636 607232 312688 607238
rect 312636 607174 312688 607180
rect 312648 555558 312676 607174
rect 313936 561134 313964 635122
rect 314016 635044 314068 635050
rect 314016 634986 314068 634992
rect 314028 568206 314056 634986
rect 314200 633956 314252 633962
rect 314200 633898 314252 633904
rect 314108 633684 314160 633690
rect 314108 633626 314160 633632
rect 314016 568200 314068 568206
rect 314016 568142 314068 568148
rect 314120 567730 314148 633626
rect 314108 567724 314160 567730
rect 314108 567666 314160 567672
rect 314212 567662 314240 633898
rect 316684 616888 316736 616894
rect 316684 616830 316736 616836
rect 314200 567656 314252 567662
rect 314200 567598 314252 567604
rect 313924 561128 313976 561134
rect 313924 561070 313976 561076
rect 312636 555552 312688 555558
rect 312636 555494 312688 555500
rect 312544 554192 312596 554198
rect 312544 554134 312596 554140
rect 311256 552968 311308 552974
rect 311256 552910 311308 552916
rect 313924 552356 313976 552362
rect 313924 552298 313976 552304
rect 307024 551268 307076 551274
rect 307024 551210 307076 551216
rect 305644 520872 305696 520878
rect 305644 520814 305696 520820
rect 307036 519926 307064 551210
rect 307024 519920 307076 519926
rect 307024 519862 307076 519868
rect 304448 519444 304500 519450
rect 304448 519386 304500 519392
rect 302976 518220 303028 518226
rect 302976 518162 303028 518168
rect 313936 517478 313964 552298
rect 313924 517472 313976 517478
rect 313924 517414 313976 517420
rect 302698 510504 302754 510513
rect 302698 510439 302754 510448
rect 302238 495544 302294 495553
rect 302238 495479 302240 495488
rect 302292 495479 302294 495488
rect 302240 495450 302292 495456
rect 59372 488022 60214 488050
rect 60598 488022 60688 488050
rect 56416 485784 56468 485790
rect 56416 485726 56468 485732
rect 56324 485444 56376 485450
rect 56324 485386 56376 485392
rect 54668 485308 54720 485314
rect 54668 485250 54720 485256
rect 53656 484968 53708 484974
rect 53656 484910 53708 484916
rect 53288 484832 53340 484838
rect 53288 484774 53340 484780
rect 53300 484537 53328 484774
rect 53668 484537 53696 484910
rect 53286 484528 53342 484537
rect 53286 484463 53342 484472
rect 53654 484528 53710 484537
rect 53654 484463 53710 484472
rect 54576 482180 54628 482186
rect 54576 482122 54628 482128
rect 54484 479460 54536 479466
rect 54484 479402 54536 479408
rect 53288 479392 53340 479398
rect 53288 479334 53340 479340
rect 53196 474428 53248 474434
rect 53196 474370 53248 474376
rect 53104 471436 53156 471442
rect 53104 471378 53156 471384
rect 53012 471300 53064 471306
rect 53012 471242 53064 471248
rect 52920 464500 52972 464506
rect 52920 464442 52972 464448
rect 52368 389156 52420 389162
rect 52368 389098 52420 389104
rect 52366 388512 52422 388521
rect 52366 388447 52422 388456
rect 52276 59424 52328 59430
rect 52276 59366 52328 59372
rect 52380 57662 52408 388447
rect 52932 380730 52960 464442
rect 52920 380724 52972 380730
rect 52920 380666 52972 380672
rect 52920 282396 52972 282402
rect 52920 282338 52972 282344
rect 52458 272776 52514 272785
rect 52458 272711 52514 272720
rect 52472 271726 52500 272711
rect 52736 272060 52788 272066
rect 52736 272002 52788 272008
rect 52460 271720 52512 271726
rect 52460 271662 52512 271668
rect 52748 270230 52776 272002
rect 52828 271720 52880 271726
rect 52828 271662 52880 271668
rect 52736 270224 52788 270230
rect 52736 270166 52788 270172
rect 52840 267734 52868 271662
rect 52932 271250 52960 282338
rect 53024 277394 53052 471242
rect 53116 282282 53144 471378
rect 53208 282402 53236 474370
rect 53196 282396 53248 282402
rect 53196 282338 53248 282344
rect 53116 282254 53236 282282
rect 53024 277366 53144 277394
rect 53010 271824 53066 271833
rect 53010 271759 53066 271768
rect 52920 271244 52972 271250
rect 52920 271186 52972 271192
rect 52840 267706 52960 267734
rect 52932 148646 52960 267706
rect 52920 148640 52972 148646
rect 52920 148582 52972 148588
rect 53024 58682 53052 271759
rect 53116 271522 53144 277366
rect 53104 271516 53156 271522
rect 53104 271458 53156 271464
rect 53208 271386 53236 282254
rect 53300 272066 53328 479334
rect 53380 479324 53432 479330
rect 53380 479266 53432 479272
rect 53288 272060 53340 272066
rect 53288 272002 53340 272008
rect 53392 271810 53420 479266
rect 53564 471912 53616 471918
rect 53564 471854 53616 471860
rect 53472 468716 53524 468722
rect 53472 468658 53524 468664
rect 53300 271782 53420 271810
rect 53196 271380 53248 271386
rect 53196 271322 53248 271328
rect 53300 270586 53328 271782
rect 53208 270558 53328 270586
rect 53208 270434 53236 270558
rect 53286 270464 53342 270473
rect 53196 270428 53248 270434
rect 53286 270399 53342 270408
rect 53196 270370 53248 270376
rect 53104 148368 53156 148374
rect 53104 148310 53156 148316
rect 53012 58676 53064 58682
rect 53012 58618 53064 58624
rect 52368 57656 52420 57662
rect 52368 57598 52420 57604
rect 53116 56506 53144 148310
rect 53208 146198 53236 270370
rect 53196 146192 53248 146198
rect 53196 146134 53248 146140
rect 53104 56500 53156 56506
rect 53104 56442 53156 56448
rect 52184 55072 52236 55078
rect 52184 55014 52236 55020
rect 53208 54874 53236 146134
rect 53300 144770 53328 270399
rect 53484 164830 53512 468658
rect 53576 166802 53604 471854
rect 53656 471708 53708 471714
rect 53656 471650 53708 471656
rect 53564 166796 53616 166802
rect 53564 166738 53616 166744
rect 53472 164824 53524 164830
rect 53472 164766 53524 164772
rect 53668 163946 53696 471650
rect 54392 466200 54444 466206
rect 54392 466142 54444 466148
rect 54300 466064 54352 466070
rect 54300 466006 54352 466012
rect 53748 465792 53800 465798
rect 53748 465734 53800 465740
rect 53656 163940 53708 163946
rect 53656 163882 53708 163888
rect 53656 163600 53708 163606
rect 53656 163542 53708 163548
rect 53472 148776 53524 148782
rect 53472 148718 53524 148724
rect 53288 144764 53340 144770
rect 53288 144706 53340 144712
rect 53484 55894 53512 148718
rect 53564 148436 53616 148442
rect 53564 148378 53616 148384
rect 53472 55888 53524 55894
rect 53472 55830 53524 55836
rect 53576 55146 53604 148378
rect 53668 56370 53696 163542
rect 53760 57730 53788 465734
rect 54312 378010 54340 466006
rect 54404 378078 54432 466142
rect 54392 378072 54444 378078
rect 54392 378014 54444 378020
rect 54300 378004 54352 378010
rect 54300 377946 54352 377952
rect 54390 375456 54446 375465
rect 54390 375391 54446 375400
rect 54300 358080 54352 358086
rect 54300 358022 54352 358028
rect 54206 282296 54262 282305
rect 54206 282231 54262 282240
rect 53840 271448 53892 271454
rect 53840 271390 53892 271396
rect 53852 271153 53880 271390
rect 53838 271144 53894 271153
rect 53838 271079 53894 271088
rect 53840 251864 53892 251870
rect 53840 251806 53892 251812
rect 53852 251122 53880 251806
rect 53840 251116 53892 251122
rect 53840 251058 53892 251064
rect 53748 57724 53800 57730
rect 53748 57666 53800 57672
rect 54220 57594 54248 282231
rect 54312 271726 54340 358022
rect 54404 282198 54432 375391
rect 54392 282192 54444 282198
rect 54392 282134 54444 282140
rect 54300 271720 54352 271726
rect 54300 271662 54352 271668
rect 54390 271144 54446 271153
rect 54390 271079 54446 271088
rect 54300 251116 54352 251122
rect 54300 251058 54352 251064
rect 54312 165646 54340 251058
rect 54404 166258 54432 271079
rect 54496 270026 54524 479402
rect 54588 270978 54616 482122
rect 54680 271590 54708 485250
rect 56232 485104 56284 485110
rect 56232 485046 56284 485052
rect 55772 477284 55824 477290
rect 55772 477226 55824 477232
rect 54760 474496 54812 474502
rect 54760 474438 54812 474444
rect 54668 271584 54720 271590
rect 54668 271526 54720 271532
rect 54772 271454 54800 474438
rect 55126 471608 55182 471617
rect 55126 471543 55182 471552
rect 54944 469056 54996 469062
rect 54944 468998 54996 469004
rect 54852 468852 54904 468858
rect 54852 468794 54904 468800
rect 54760 271448 54812 271454
rect 54760 271390 54812 271396
rect 54576 270972 54628 270978
rect 54576 270914 54628 270920
rect 54576 270224 54628 270230
rect 54576 270166 54628 270172
rect 54484 270020 54536 270026
rect 54484 269962 54536 269968
rect 54484 252000 54536 252006
rect 54484 251942 54536 251948
rect 54392 166252 54444 166258
rect 54392 166194 54444 166200
rect 54300 165640 54352 165646
rect 54300 165582 54352 165588
rect 54208 57588 54260 57594
rect 54208 57530 54260 57536
rect 54312 56574 54340 165582
rect 54496 145897 54524 251942
rect 54482 145888 54538 145897
rect 54588 145858 54616 270166
rect 54668 269748 54720 269754
rect 54668 269690 54720 269696
rect 54482 145823 54538 145832
rect 54576 145852 54628 145858
rect 54576 145794 54628 145800
rect 54392 145648 54444 145654
rect 54392 145590 54444 145596
rect 54574 145616 54630 145625
rect 54404 59702 54432 145590
rect 54574 145551 54630 145560
rect 54484 145444 54536 145450
rect 54484 145386 54536 145392
rect 54496 59770 54524 145386
rect 54484 59764 54536 59770
rect 54484 59706 54536 59712
rect 54392 59696 54444 59702
rect 54392 59638 54444 59644
rect 54588 59566 54616 145551
rect 54680 144906 54708 269690
rect 54864 165374 54892 468794
rect 54852 165368 54904 165374
rect 54852 165310 54904 165316
rect 54956 164966 54984 468998
rect 55036 468920 55088 468926
rect 55036 468862 55088 468868
rect 55048 165170 55076 468862
rect 55140 165442 55168 471543
rect 55680 466336 55732 466342
rect 55680 466278 55732 466284
rect 55692 465225 55720 466278
rect 55678 465216 55734 465225
rect 55678 465151 55734 465160
rect 55680 418260 55732 418266
rect 55680 418202 55732 418208
rect 55692 417466 55720 418202
rect 55784 418198 55812 477226
rect 56138 471336 56194 471345
rect 56138 471271 56194 471280
rect 56048 468988 56100 468994
rect 56048 468930 56100 468936
rect 55864 464568 55916 464574
rect 55864 464510 55916 464516
rect 55772 418192 55824 418198
rect 55772 418134 55824 418140
rect 55692 417438 55812 417466
rect 55680 415404 55732 415410
rect 55680 415346 55732 415352
rect 55692 381070 55720 415346
rect 55680 381064 55732 381070
rect 55680 381006 55732 381012
rect 55784 378894 55812 417438
rect 55876 380934 55904 464510
rect 55956 464364 56008 464370
rect 55956 464306 56008 464312
rect 55864 380928 55916 380934
rect 55864 380870 55916 380876
rect 55864 380724 55916 380730
rect 55864 380666 55916 380672
rect 55772 378888 55824 378894
rect 55772 378830 55824 378836
rect 55876 282742 55904 380666
rect 55968 379302 55996 464306
rect 55956 379296 56008 379302
rect 55956 379238 56008 379244
rect 55864 282736 55916 282742
rect 55864 282678 55916 282684
rect 55956 270020 56008 270026
rect 55956 269962 56008 269968
rect 55128 165436 55180 165442
rect 55128 165378 55180 165384
rect 55036 165164 55088 165170
rect 55036 165106 55088 165112
rect 54944 164960 54996 164966
rect 54944 164902 54996 164908
rect 55036 163736 55088 163742
rect 55036 163678 55088 163684
rect 54944 148844 54996 148850
rect 54944 148786 54996 148792
rect 54852 145852 54904 145858
rect 54852 145794 54904 145800
rect 54760 145376 54812 145382
rect 54760 145318 54812 145324
rect 54668 144900 54720 144906
rect 54668 144842 54720 144848
rect 54576 59560 54628 59566
rect 54576 59502 54628 59508
rect 54772 57186 54800 145318
rect 54760 57180 54812 57186
rect 54760 57122 54812 57128
rect 54300 56568 54352 56574
rect 54300 56510 54352 56516
rect 53656 56364 53708 56370
rect 53656 56306 53708 56312
rect 54864 56098 54892 145794
rect 54852 56092 54904 56098
rect 54852 56034 54904 56040
rect 53564 55140 53616 55146
rect 53564 55082 53616 55088
rect 53196 54868 53248 54874
rect 53196 54810 53248 54816
rect 54956 54670 54984 148786
rect 55048 59090 55076 163678
rect 55968 151814 55996 269962
rect 56060 165102 56088 468930
rect 56152 165510 56180 471271
rect 56244 166598 56272 485046
rect 56232 166592 56284 166598
rect 56232 166534 56284 166540
rect 56140 165504 56192 165510
rect 56140 165446 56192 165452
rect 56336 165238 56364 485386
rect 56324 165232 56376 165238
rect 56324 165174 56376 165180
rect 56048 165096 56100 165102
rect 56048 165038 56100 165044
rect 56428 164694 56456 485726
rect 56508 485580 56560 485586
rect 56508 485522 56560 485528
rect 56520 165306 56548 485522
rect 58624 485036 58676 485042
rect 58624 484978 58676 484984
rect 56784 483676 56836 483682
rect 56784 483618 56836 483624
rect 56796 307737 56824 483618
rect 57244 482316 57296 482322
rect 57244 482258 57296 482264
rect 57152 476740 57204 476746
rect 57152 476682 57204 476688
rect 57060 464432 57112 464438
rect 57060 464374 57112 464380
rect 56876 418192 56928 418198
rect 56876 418134 56928 418140
rect 56888 412634 56916 418134
rect 56968 418124 57020 418130
rect 56968 418066 57020 418072
rect 56980 417217 57008 418066
rect 56966 417208 57022 417217
rect 56966 417143 57022 417152
rect 57072 415410 57100 464374
rect 57164 418266 57192 476682
rect 57152 418260 57204 418266
rect 57152 418202 57204 418208
rect 57060 415404 57112 415410
rect 57060 415346 57112 415352
rect 57152 415404 57204 415410
rect 57152 415346 57204 415352
rect 56888 412606 57008 412634
rect 56980 386374 57008 412606
rect 57060 391944 57112 391950
rect 57060 391886 57112 391892
rect 57072 391513 57100 391886
rect 57058 391504 57114 391513
rect 57058 391439 57114 391448
rect 57060 389088 57112 389094
rect 57058 389056 57060 389065
rect 57112 389056 57114 389065
rect 57058 388991 57114 389000
rect 56968 386368 57020 386374
rect 56968 386310 57020 386316
rect 57164 378962 57192 415346
rect 57256 413982 57284 482258
rect 57796 481024 57848 481030
rect 57796 480966 57848 480972
rect 57336 477352 57388 477358
rect 57336 477294 57388 477300
rect 57244 413976 57296 413982
rect 57244 413918 57296 413924
rect 57244 389156 57296 389162
rect 57244 389098 57296 389104
rect 57152 378956 57204 378962
rect 57152 378898 57204 378904
rect 57152 357876 57204 357882
rect 57152 357818 57204 357824
rect 56874 309088 56930 309097
rect 56874 309023 56930 309032
rect 56888 307873 56916 309023
rect 56874 307864 56930 307873
rect 56874 307799 56930 307808
rect 56782 307728 56838 307737
rect 56782 307663 56838 307672
rect 56782 203552 56838 203561
rect 56782 203487 56838 203496
rect 56508 165300 56560 165306
rect 56508 165242 56560 165248
rect 56416 164688 56468 164694
rect 56416 164630 56468 164636
rect 56508 163804 56560 163810
rect 56508 163746 56560 163752
rect 55968 151786 56180 151814
rect 55864 148640 55916 148646
rect 55864 148582 55916 148588
rect 55036 59084 55088 59090
rect 55036 59026 55088 59032
rect 55876 58954 55904 148582
rect 56152 145994 56180 151786
rect 56230 146296 56286 146305
rect 56230 146231 56286 146240
rect 56140 145988 56192 145994
rect 56140 145930 56192 145936
rect 56048 144900 56100 144906
rect 56048 144842 56100 144848
rect 55956 144696 56008 144702
rect 55956 144638 56008 144644
rect 55864 58948 55916 58954
rect 55864 58890 55916 58896
rect 55968 57390 55996 144638
rect 56060 59362 56088 144842
rect 56152 144514 56180 145930
rect 56244 144634 56272 146231
rect 56322 145752 56378 145761
rect 56322 145687 56378 145696
rect 56416 145716 56468 145722
rect 56336 144702 56364 145687
rect 56416 145658 56468 145664
rect 56428 144906 56456 145658
rect 56416 144900 56468 144906
rect 56416 144842 56468 144848
rect 56324 144696 56376 144702
rect 56324 144638 56376 144644
rect 56232 144628 56284 144634
rect 56232 144570 56284 144576
rect 56152 144486 56456 144514
rect 56324 144424 56376 144430
rect 56324 144366 56376 144372
rect 56048 59356 56100 59362
rect 56048 59298 56100 59304
rect 56336 59022 56364 144366
rect 56324 59016 56376 59022
rect 56324 58958 56376 58964
rect 55956 57384 56008 57390
rect 55956 57326 56008 57332
rect 56428 56166 56456 144486
rect 56520 59158 56548 163746
rect 56796 96529 56824 203487
rect 56888 201385 56916 307799
rect 57060 300824 57112 300830
rect 57060 300766 57112 300772
rect 56968 252476 57020 252482
rect 56968 252418 57020 252424
rect 56874 201376 56930 201385
rect 56874 201311 56930 201320
rect 56980 164014 57008 252418
rect 57072 195265 57100 300766
rect 57164 271658 57192 357818
rect 57256 282577 57284 389098
rect 57348 387802 57376 477294
rect 57428 474360 57480 474366
rect 57428 474302 57480 474308
rect 57336 387796 57388 387802
rect 57336 387738 57388 387744
rect 57440 381682 57468 474302
rect 57704 474156 57756 474162
rect 57704 474098 57756 474104
rect 57520 471368 57572 471374
rect 57520 471310 57572 471316
rect 57532 389434 57560 471310
rect 57612 469872 57664 469878
rect 57612 469814 57664 469820
rect 57520 389428 57572 389434
rect 57520 389370 57572 389376
rect 57518 389328 57574 389337
rect 57518 389263 57574 389272
rect 57532 389162 57560 389263
rect 57520 389156 57572 389162
rect 57520 389098 57572 389104
rect 57520 389020 57572 389026
rect 57520 388962 57572 388968
rect 57428 381676 57480 381682
rect 57428 381618 57480 381624
rect 57532 311137 57560 388962
rect 57518 311128 57574 311137
rect 57518 311063 57574 311072
rect 57334 310448 57390 310457
rect 57334 310383 57390 310392
rect 57242 282568 57298 282577
rect 57242 282503 57298 282512
rect 57152 271652 57204 271658
rect 57152 271594 57204 271600
rect 57244 269884 57296 269890
rect 57244 269826 57296 269832
rect 57256 268977 57284 269826
rect 57242 268968 57298 268977
rect 57242 268903 57298 268912
rect 57150 204232 57206 204241
rect 57150 204167 57206 204176
rect 57058 195256 57114 195265
rect 57058 195191 57114 195200
rect 56968 164008 57020 164014
rect 56968 163950 57020 163956
rect 57060 163872 57112 163878
rect 57060 163814 57112 163820
rect 56968 146260 57020 146266
rect 56968 146202 57020 146208
rect 56782 96520 56838 96529
rect 56782 96455 56838 96464
rect 56508 59152 56560 59158
rect 56508 59094 56560 59100
rect 56416 56160 56468 56166
rect 56416 56102 56468 56108
rect 56980 54942 57008 146202
rect 57072 59226 57100 163814
rect 57164 97481 57192 204167
rect 57256 146266 57284 268903
rect 57348 203561 57376 310383
rect 57426 301608 57482 301617
rect 57426 301543 57482 301552
rect 57440 300830 57468 301543
rect 57428 300824 57480 300830
rect 57428 300766 57480 300772
rect 57428 300688 57480 300694
rect 57428 300630 57480 300636
rect 57334 203552 57390 203561
rect 57334 203487 57390 203496
rect 57334 198792 57390 198801
rect 57334 198727 57390 198736
rect 57244 146260 57296 146266
rect 57244 146202 57296 146208
rect 57150 97472 57206 97481
rect 57150 97407 57206 97416
rect 57348 93401 57376 198727
rect 57440 196353 57468 300630
rect 57532 204241 57560 311063
rect 57624 306374 57652 469814
rect 57716 309097 57744 474098
rect 57808 310457 57836 480966
rect 58440 476672 58492 476678
rect 58440 476614 58492 476620
rect 57886 417344 57942 417353
rect 57886 417279 57942 417288
rect 57900 416838 57928 417279
rect 57888 416832 57940 416838
rect 57888 416774 57940 416780
rect 58452 415410 58480 476614
rect 58532 476604 58584 476610
rect 58532 476546 58584 476552
rect 58440 415404 58492 415410
rect 58440 415346 58492 415352
rect 57886 414216 57942 414225
rect 57886 414151 57942 414160
rect 57900 414050 57928 414151
rect 57888 414044 57940 414050
rect 57888 413986 57940 413992
rect 58440 413976 58492 413982
rect 58440 413918 58492 413924
rect 57886 413264 57942 413273
rect 57886 413199 57942 413208
rect 57900 412690 57928 413199
rect 57888 412684 57940 412690
rect 57888 412626 57940 412632
rect 57886 411496 57942 411505
rect 57886 411431 57942 411440
rect 57900 411330 57928 411431
rect 57888 411324 57940 411330
rect 57888 411266 57940 411272
rect 57886 410408 57942 410417
rect 57886 410343 57942 410352
rect 57900 409902 57928 410343
rect 57888 409896 57940 409902
rect 57888 409838 57940 409844
rect 57886 408640 57942 408649
rect 57886 408575 57942 408584
rect 57900 408542 57928 408575
rect 57888 408536 57940 408542
rect 57888 408478 57940 408484
rect 57888 387184 57940 387190
rect 57888 387126 57940 387132
rect 57900 380458 57928 387126
rect 57888 380452 57940 380458
rect 57888 380394 57940 380400
rect 58452 380322 58480 413918
rect 58544 387734 58572 476546
rect 58636 388521 58664 484978
rect 59176 484900 59228 484906
rect 59176 484842 59228 484848
rect 58808 482112 58860 482118
rect 58808 482054 58860 482060
rect 58716 472864 58768 472870
rect 58716 472806 58768 472812
rect 58622 388512 58678 388521
rect 58622 388447 58678 388456
rect 58624 387796 58676 387802
rect 58624 387738 58676 387744
rect 58532 387728 58584 387734
rect 58532 387670 58584 387676
rect 58440 380316 58492 380322
rect 58440 380258 58492 380264
rect 58636 380254 58664 387738
rect 58624 380248 58676 380254
rect 58624 380190 58676 380196
rect 58532 356244 58584 356250
rect 58532 356186 58584 356192
rect 57794 310448 57850 310457
rect 57794 310383 57850 310392
rect 57702 309088 57758 309097
rect 57702 309023 57758 309032
rect 57794 307728 57850 307737
rect 57794 307663 57850 307672
rect 57808 306785 57836 307663
rect 57794 306776 57850 306785
rect 57794 306711 57850 306720
rect 57624 306346 57744 306374
rect 57716 305017 57744 306346
rect 57702 305008 57758 305017
rect 57702 304943 57758 304952
rect 57610 303648 57666 303657
rect 57610 303583 57612 303592
rect 57664 303583 57666 303592
rect 57612 303554 57664 303560
rect 57624 300694 57652 303554
rect 57612 300688 57664 300694
rect 57612 300630 57664 300636
rect 57518 204232 57574 204241
rect 57518 204167 57574 204176
rect 57610 201376 57666 201385
rect 57610 201311 57666 201320
rect 57426 196344 57482 196353
rect 57426 196279 57482 196288
rect 57334 93392 57390 93401
rect 57334 93327 57390 93336
rect 57440 90545 57468 196279
rect 57520 164144 57572 164150
rect 57518 164112 57520 164121
rect 57572 164112 57574 164121
rect 57518 164047 57574 164056
rect 57624 93809 57652 201311
rect 57716 198234 57744 304943
rect 57808 199889 57836 306711
rect 58440 282736 58492 282742
rect 58440 282678 58492 282684
rect 57886 282568 57942 282577
rect 57886 282503 57942 282512
rect 57794 199880 57850 199889
rect 57794 199815 57850 199824
rect 57808 198801 57836 199815
rect 57794 198792 57850 198801
rect 57794 198727 57850 198736
rect 57716 198206 57836 198234
rect 57808 198121 57836 198206
rect 57794 198112 57850 198121
rect 57794 198047 57850 198056
rect 57702 195256 57758 195265
rect 57702 195191 57758 195200
rect 57610 93800 57666 93809
rect 57610 93735 57666 93744
rect 57426 90536 57482 90545
rect 57426 90471 57482 90480
rect 57716 88233 57744 195191
rect 57808 91089 57836 198047
rect 57900 175817 57928 282503
rect 58452 272270 58480 282678
rect 58544 281518 58572 356186
rect 58624 356040 58676 356046
rect 58624 355982 58676 355988
rect 58532 281512 58584 281518
rect 58532 281454 58584 281460
rect 58636 272406 58664 355982
rect 58728 284209 58756 472806
rect 58714 284200 58770 284209
rect 58714 284135 58770 284144
rect 58716 282192 58768 282198
rect 58716 282134 58768 282140
rect 58624 272400 58676 272406
rect 58624 272342 58676 272348
rect 58440 272264 58492 272270
rect 58440 272206 58492 272212
rect 58728 272202 58756 282134
rect 58820 282033 58848 482054
rect 58900 471504 58952 471510
rect 58900 471446 58952 471452
rect 58806 282024 58862 282033
rect 58806 281959 58862 281968
rect 58716 272196 58768 272202
rect 58716 272138 58768 272144
rect 58624 270156 58676 270162
rect 58624 270098 58676 270104
rect 58636 269074 58664 270098
rect 58624 269068 58676 269074
rect 58624 269010 58676 269016
rect 58532 251932 58584 251938
rect 58532 251874 58584 251880
rect 58544 251190 58572 251874
rect 58532 251184 58584 251190
rect 58532 251126 58584 251132
rect 57886 175808 57942 175817
rect 57886 175743 57942 175752
rect 57794 91080 57850 91089
rect 57794 91015 57850 91024
rect 57702 88224 57758 88233
rect 57702 88159 57758 88168
rect 57612 70372 57664 70378
rect 57612 70314 57664 70320
rect 57624 70145 57652 70314
rect 57610 70136 57666 70145
rect 57610 70071 57666 70080
rect 57900 68921 57928 175743
rect 58544 164218 58572 251126
rect 58532 164212 58584 164218
rect 58532 164154 58584 164160
rect 58636 146130 58664 269010
rect 58808 252544 58860 252550
rect 58808 252486 58860 252492
rect 58716 251660 58768 251666
rect 58716 251602 58768 251608
rect 58728 149054 58756 251602
rect 58716 149048 58768 149054
rect 58716 148990 58768 148996
rect 58728 147801 58756 148990
rect 58714 147792 58770 147801
rect 58714 147727 58770 147736
rect 58820 146305 58848 252486
rect 58912 177585 58940 471446
rect 59084 464704 59136 464710
rect 59084 464646 59136 464652
rect 58992 464636 59044 464642
rect 58992 464578 59044 464584
rect 58898 177576 58954 177585
rect 58898 177511 58954 177520
rect 59004 166394 59032 464578
rect 59096 166666 59124 464646
rect 59084 166660 59136 166666
rect 59084 166602 59136 166608
rect 59188 166462 59216 484842
rect 59372 474026 59400 488022
rect 59912 485648 59964 485654
rect 59912 485590 59964 485596
rect 59636 480072 59688 480078
rect 59636 480014 59688 480020
rect 59360 474020 59412 474026
rect 59360 473962 59412 473968
rect 59268 466132 59320 466138
rect 59268 466074 59320 466080
rect 59176 166456 59228 166462
rect 59176 166398 59228 166404
rect 58992 166388 59044 166394
rect 58992 166330 59044 166336
rect 59176 148504 59228 148510
rect 59176 148446 59228 148452
rect 59188 147626 59216 148446
rect 58900 147620 58952 147626
rect 58900 147562 58952 147568
rect 59176 147620 59228 147626
rect 59176 147562 59228 147568
rect 58806 146296 58862 146305
rect 58806 146231 58862 146240
rect 58624 146124 58676 146130
rect 58624 146066 58676 146072
rect 58716 145784 58768 145790
rect 58716 145726 58768 145732
rect 58624 145580 58676 145586
rect 58624 145522 58676 145528
rect 58636 144770 58664 145522
rect 58728 144838 58756 145726
rect 58716 144832 58768 144838
rect 58716 144774 58768 144780
rect 58624 144764 58676 144770
rect 58624 144706 58676 144712
rect 57886 68912 57942 68921
rect 57886 68847 57942 68856
rect 57060 59220 57112 59226
rect 57060 59162 57112 59168
rect 57900 57934 57928 68847
rect 57888 57928 57940 57934
rect 57888 57870 57940 57876
rect 57900 57526 57928 57870
rect 57244 57520 57296 57526
rect 57244 57462 57296 57468
rect 57888 57520 57940 57526
rect 57888 57462 57940 57468
rect 56968 54936 57020 54942
rect 56968 54878 57020 54884
rect 54944 54664 54996 54670
rect 54944 54606 54996 54612
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 10324 20664 10376 20670
rect 10324 20606 10376 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 57256 3466 57284 57462
rect 58636 56234 58664 144706
rect 58624 56228 58676 56234
rect 58624 56170 58676 56176
rect 58728 55962 58756 144774
rect 58912 59498 58940 147562
rect 59084 146260 59136 146266
rect 59084 146202 59136 146208
rect 58990 145888 59046 145897
rect 58990 145823 59046 145832
rect 59004 59634 59032 145823
rect 58992 59628 59044 59634
rect 58992 59570 59044 59576
rect 58900 59492 58952 59498
rect 58900 59434 58952 59440
rect 58716 55956 58768 55962
rect 58716 55898 58768 55904
rect 59096 54806 59124 146202
rect 59176 146124 59228 146130
rect 59176 146066 59228 146072
rect 59188 145926 59216 146066
rect 59176 145920 59228 145926
rect 59176 145862 59228 145868
rect 59084 54800 59136 54806
rect 59084 54742 59136 54748
rect 59188 54738 59216 145862
rect 59280 57322 59308 466074
rect 59360 387728 59412 387734
rect 59360 387670 59412 387676
rect 59372 356250 59400 387670
rect 59544 381676 59596 381682
rect 59544 381618 59596 381624
rect 59452 381064 59504 381070
rect 59452 381006 59504 381012
rect 59360 356244 59412 356250
rect 59360 356186 59412 356192
rect 59464 356046 59492 381006
rect 59556 357882 59584 381618
rect 59648 379438 59676 480014
rect 59728 477488 59780 477494
rect 59728 477430 59780 477436
rect 59740 387190 59768 477430
rect 59818 471744 59874 471753
rect 59818 471679 59874 471688
rect 59728 387184 59780 387190
rect 59728 387126 59780 387132
rect 59728 386368 59780 386374
rect 59728 386310 59780 386316
rect 59740 380526 59768 386310
rect 59728 380520 59780 380526
rect 59728 380462 59780 380468
rect 59636 379432 59688 379438
rect 59636 379374 59688 379380
rect 59544 357876 59596 357882
rect 59544 357818 59596 357824
rect 59452 356040 59504 356046
rect 59452 355982 59504 355988
rect 59728 281512 59780 281518
rect 59728 281454 59780 281460
rect 59450 272640 59506 272649
rect 59450 272575 59506 272584
rect 59464 272406 59492 272575
rect 59452 272400 59504 272406
rect 59452 272342 59504 272348
rect 59360 270088 59412 270094
rect 59360 270030 59412 270036
rect 59372 269113 59400 270030
rect 59358 269104 59414 269113
rect 59358 269039 59414 269048
rect 59372 146266 59400 269039
rect 59464 175953 59492 272342
rect 59740 270298 59768 281454
rect 59728 270292 59780 270298
rect 59728 270234 59780 270240
rect 59450 175944 59506 175953
rect 59450 175879 59506 175888
rect 59832 165578 59860 471679
rect 59924 166530 59952 485590
rect 60660 483750 60688 488022
rect 60740 484152 60792 484158
rect 60740 484094 60792 484100
rect 60648 483744 60700 483750
rect 60648 483686 60700 483692
rect 60752 465866 60780 484094
rect 60832 484016 60884 484022
rect 60832 483958 60884 483964
rect 60844 466002 60872 483958
rect 61028 475386 61056 488036
rect 61120 488022 61502 488050
rect 61672 488022 61962 488050
rect 62224 488022 62330 488050
rect 62408 488022 62790 488050
rect 62960 488022 63250 488050
rect 63512 488022 63710 488050
rect 61120 484158 61148 488022
rect 61108 484152 61160 484158
rect 61108 484094 61160 484100
rect 61672 484022 61700 488022
rect 62120 484152 62172 484158
rect 62120 484094 62172 484100
rect 61660 484016 61712 484022
rect 61660 483958 61712 483964
rect 61016 475380 61068 475386
rect 61016 475322 61068 475328
rect 62132 466206 62160 484094
rect 62224 478145 62252 488022
rect 62408 479534 62436 488022
rect 62960 484158 62988 488022
rect 62948 484152 63000 484158
rect 62948 484094 63000 484100
rect 62396 479528 62448 479534
rect 62396 479470 62448 479476
rect 62210 478136 62266 478145
rect 62210 478071 62266 478080
rect 62120 466200 62172 466206
rect 62120 466142 62172 466148
rect 63512 466070 63540 488022
rect 64156 485382 64184 488036
rect 64248 488022 64538 488050
rect 64144 485376 64196 485382
rect 64144 485318 64196 485324
rect 64248 470594 64276 488022
rect 64880 484152 64932 484158
rect 64880 484094 64932 484100
rect 64892 471170 64920 484094
rect 64880 471164 64932 471170
rect 64880 471106 64932 471112
rect 64984 471102 65012 488036
rect 65076 488022 65458 488050
rect 65536 488022 65918 488050
rect 65076 471238 65104 488022
rect 65536 484158 65564 488022
rect 65524 484152 65576 484158
rect 65524 484094 65576 484100
rect 66364 482905 66392 488036
rect 66456 488022 66746 488050
rect 66824 488022 67206 488050
rect 66350 482896 66406 482905
rect 66350 482831 66406 482840
rect 66456 482746 66484 488022
rect 66272 482718 66484 482746
rect 65064 471232 65116 471238
rect 65064 471174 65116 471180
rect 64972 471096 65024 471102
rect 64972 471038 65024 471044
rect 63604 470566 64276 470594
rect 63604 468450 63632 470566
rect 63592 468444 63644 468450
rect 63592 468386 63644 468392
rect 66272 466449 66300 482718
rect 66824 470594 66852 488022
rect 66364 470566 66852 470594
rect 66258 466440 66314 466449
rect 66258 466375 66314 466384
rect 63500 466064 63552 466070
rect 63500 466006 63552 466012
rect 60832 465996 60884 466002
rect 60832 465938 60884 465944
rect 60740 465860 60792 465866
rect 60740 465802 60792 465808
rect 66364 465730 66392 470566
rect 67652 466138 67680 488036
rect 67836 488022 68126 488050
rect 68204 488022 68494 488050
rect 67732 484152 67784 484158
rect 67732 484094 67784 484100
rect 67744 469169 67772 484094
rect 67836 469849 67864 488022
rect 68204 484158 68232 488022
rect 68940 484945 68968 488036
rect 69124 488022 69414 488050
rect 69584 488022 69874 488050
rect 69952 488022 70334 488050
rect 70596 488022 70702 488050
rect 70872 488022 71162 488050
rect 71240 488022 71622 488050
rect 71792 488022 72082 488050
rect 68926 484936 68982 484945
rect 68926 484871 68982 484880
rect 68284 484764 68336 484770
rect 68284 484706 68336 484712
rect 68192 484152 68244 484158
rect 68192 484094 68244 484100
rect 67822 469840 67878 469849
rect 67822 469775 67878 469784
rect 68296 469198 68324 484706
rect 69020 484152 69072 484158
rect 69020 484094 69072 484100
rect 68284 469192 68336 469198
rect 67730 469160 67786 469169
rect 68284 469134 68336 469140
rect 67730 469095 67786 469104
rect 67640 466132 67692 466138
rect 67640 466074 67692 466080
rect 69032 465905 69060 484094
rect 69018 465896 69074 465905
rect 69018 465831 69074 465840
rect 66352 465724 66404 465730
rect 66352 465666 66404 465672
rect 69124 465633 69152 488022
rect 69584 484158 69612 488022
rect 69664 485512 69716 485518
rect 69664 485454 69716 485460
rect 69676 484906 69704 485454
rect 69664 484900 69716 484906
rect 69664 484842 69716 484848
rect 69572 484152 69624 484158
rect 69572 484094 69624 484100
rect 69952 470594 69980 488022
rect 70400 480888 70452 480894
rect 70400 480830 70452 480836
rect 69216 470566 69980 470594
rect 69216 469033 69244 470566
rect 69202 469024 69258 469033
rect 69202 468959 69258 468968
rect 70412 465934 70440 480830
rect 70492 480820 70544 480826
rect 70492 480762 70544 480768
rect 70504 467362 70532 480762
rect 70596 469130 70624 488022
rect 70872 480894 70900 488022
rect 70860 480888 70912 480894
rect 70860 480830 70912 480836
rect 71240 480826 71268 488022
rect 71228 480820 71280 480826
rect 71228 480762 71280 480768
rect 70584 469124 70636 469130
rect 70584 469066 70636 469072
rect 70492 467356 70544 467362
rect 70492 467298 70544 467304
rect 71792 466313 71820 488022
rect 72528 485761 72556 488036
rect 72620 488022 72910 488050
rect 73172 488022 73370 488050
rect 72514 485752 72570 485761
rect 72514 485687 72570 485696
rect 72620 485466 72648 488022
rect 71884 485438 72648 485466
rect 71884 467129 71912 485438
rect 72424 485376 72476 485382
rect 72424 485318 72476 485324
rect 71870 467120 71926 467129
rect 71870 467055 71926 467064
rect 71778 466304 71834 466313
rect 71778 466239 71834 466248
rect 70400 465928 70452 465934
rect 70400 465870 70452 465876
rect 72436 465730 72464 485318
rect 73172 467265 73200 488022
rect 73816 485625 73844 488036
rect 73896 485716 73948 485722
rect 73896 485658 73948 485664
rect 73802 485616 73858 485625
rect 73802 485551 73858 485560
rect 73908 485466 73936 485658
rect 74276 485489 74304 488036
rect 74674 488022 74764 488050
rect 73816 485438 73936 485466
rect 74262 485480 74318 485489
rect 73816 467294 73844 485438
rect 74262 485415 74318 485424
rect 74446 485480 74502 485489
rect 74446 485415 74502 485424
rect 73896 485376 73948 485382
rect 73896 485318 73948 485324
rect 73908 474570 73936 485318
rect 74460 484974 74488 485415
rect 74448 484968 74500 484974
rect 74448 484910 74500 484916
rect 74736 481098 74764 488022
rect 74828 488022 75118 488050
rect 75288 488022 75578 488050
rect 74724 481092 74776 481098
rect 74724 481034 74776 481040
rect 74828 480978 74856 488022
rect 74908 481092 74960 481098
rect 74908 481034 74960 481040
rect 74552 480950 74856 480978
rect 73896 474564 73948 474570
rect 73896 474506 73948 474512
rect 73804 467288 73856 467294
rect 73158 467256 73214 467265
rect 73804 467230 73856 467236
rect 73158 467191 73214 467200
rect 74552 466177 74580 480950
rect 74632 480888 74684 480894
rect 74632 480830 74684 480836
rect 74538 466168 74594 466177
rect 74538 466103 74594 466112
rect 74644 465769 74672 480830
rect 74920 470594 74948 481034
rect 75288 480894 75316 488022
rect 76024 485353 76052 488036
rect 76208 488022 76498 488050
rect 76576 488022 76866 488050
rect 76010 485344 76066 485353
rect 76010 485279 76066 485288
rect 75276 480888 75328 480894
rect 75276 480830 75328 480836
rect 75920 480888 75972 480894
rect 75920 480830 75972 480836
rect 74736 470566 74948 470594
rect 74736 465798 74764 470566
rect 75932 466410 75960 480830
rect 76208 470594 76236 488022
rect 76576 480894 76604 488022
rect 77312 485217 77340 488036
rect 77298 485208 77354 485217
rect 77298 485143 77354 485152
rect 77772 484702 77800 488036
rect 77864 488022 78246 488050
rect 77760 484696 77812 484702
rect 77760 484638 77812 484644
rect 76564 480888 76616 480894
rect 76564 480830 76616 480836
rect 77864 470594 77892 488022
rect 76024 470566 76236 470594
rect 77496 470566 77892 470594
rect 75920 466404 75972 466410
rect 75920 466346 75972 466352
rect 76024 466041 76052 470566
rect 77496 466342 77524 470566
rect 78692 468897 78720 488036
rect 78876 488022 79074 488050
rect 79152 488022 79534 488050
rect 78772 477692 78824 477698
rect 78772 477634 78824 477640
rect 78678 468888 78734 468897
rect 78678 468823 78734 468832
rect 78784 468761 78812 477634
rect 78770 468752 78826 468761
rect 78770 468687 78826 468696
rect 78876 468625 78904 488022
rect 79152 477698 79180 488022
rect 79980 485489 80008 488036
rect 80348 488022 80454 488050
rect 80532 488022 80822 488050
rect 79966 485480 80022 485489
rect 79966 485415 80022 485424
rect 79140 477692 79192 477698
rect 79140 477634 79192 477640
rect 80348 476114 80376 488022
rect 80532 480049 80560 488022
rect 81268 485042 81296 488036
rect 81728 485790 81756 488036
rect 81912 488022 82202 488050
rect 82280 488022 82662 488050
rect 82832 488022 83030 488050
rect 83200 488022 83490 488050
rect 83568 488022 83950 488050
rect 81716 485784 81768 485790
rect 81716 485726 81768 485732
rect 81256 485036 81308 485042
rect 81256 484978 81308 484984
rect 80704 483744 80756 483750
rect 80704 483686 80756 483692
rect 80518 480040 80574 480049
rect 80518 479975 80574 479984
rect 80256 476086 80376 476114
rect 78862 468616 78918 468625
rect 78862 468551 78918 468560
rect 80256 468489 80284 476086
rect 80242 468480 80298 468489
rect 80242 468415 80298 468424
rect 80716 467838 80744 483686
rect 81532 480888 81584 480894
rect 81532 480830 81584 480836
rect 81544 471481 81572 480830
rect 81912 471986 81940 488022
rect 82280 480894 82308 488022
rect 82268 480888 82320 480894
rect 82268 480830 82320 480836
rect 81900 471980 81952 471986
rect 81900 471922 81952 471928
rect 82832 471850 82860 488022
rect 82912 480888 82964 480894
rect 82912 480830 82964 480836
rect 82820 471844 82872 471850
rect 82820 471786 82872 471792
rect 82924 471646 82952 480830
rect 82912 471640 82964 471646
rect 82912 471582 82964 471588
rect 83200 471578 83228 488022
rect 83568 480894 83596 488022
rect 84396 484906 84424 488036
rect 84488 488022 84870 488050
rect 84948 488022 85238 488050
rect 85714 488022 85804 488050
rect 84384 484900 84436 484906
rect 84384 484842 84436 484848
rect 83556 480888 83608 480894
rect 83556 480830 83608 480836
rect 84292 480888 84344 480894
rect 84292 480830 84344 480836
rect 84304 471782 84332 480830
rect 84488 471918 84516 488022
rect 84948 480894 84976 488022
rect 85776 483014 85804 488022
rect 85684 482986 85804 483014
rect 85868 488022 86158 488050
rect 86328 488022 86618 488050
rect 84936 480888 84988 480894
rect 84936 480830 84988 480836
rect 85580 479188 85632 479194
rect 85580 479130 85632 479136
rect 84476 471912 84528 471918
rect 84476 471854 84528 471860
rect 84292 471776 84344 471782
rect 84292 471718 84344 471724
rect 83188 471572 83240 471578
rect 83188 471514 83240 471520
rect 81530 471472 81586 471481
rect 81530 471407 81586 471416
rect 85592 468790 85620 479130
rect 85684 478258 85712 482986
rect 85684 478230 85804 478258
rect 85672 478168 85724 478174
rect 85672 478110 85724 478116
rect 85684 469062 85712 478110
rect 85776 471714 85804 478230
rect 85868 478174 85896 488022
rect 86328 479194 86356 488022
rect 86960 480888 87012 480894
rect 86960 480830 87012 480836
rect 86316 479188 86368 479194
rect 86316 479130 86368 479136
rect 85856 478168 85908 478174
rect 85856 478110 85908 478116
rect 85764 471708 85816 471714
rect 85764 471650 85816 471656
rect 85672 469056 85724 469062
rect 85672 468998 85724 469004
rect 86972 468926 87000 480830
rect 86960 468920 87012 468926
rect 86960 468862 87012 468868
rect 85580 468784 85632 468790
rect 85580 468726 85632 468732
rect 87064 468722 87092 488036
rect 87156 488022 87446 488050
rect 87616 488022 87906 488050
rect 87156 468994 87184 488022
rect 87616 480894 87644 488022
rect 88352 485450 88380 488036
rect 88536 488022 88826 488050
rect 88340 485444 88392 485450
rect 88340 485386 88392 485392
rect 87604 480888 87656 480894
rect 87604 480830 87656 480836
rect 88432 480888 88484 480894
rect 88432 480830 88484 480836
rect 88444 471617 88472 480830
rect 88430 471608 88486 471617
rect 88430 471543 88486 471552
rect 87144 468988 87196 468994
rect 87144 468930 87196 468936
rect 88536 468858 88564 488022
rect 89180 485586 89208 488036
rect 89272 488022 89654 488050
rect 89824 488022 90114 488050
rect 89168 485580 89220 485586
rect 89168 485522 89220 485528
rect 89272 480894 89300 488022
rect 89260 480888 89312 480894
rect 89260 480830 89312 480836
rect 89824 471345 89852 488022
rect 90560 485110 90588 488036
rect 90744 488022 91034 488050
rect 90548 485104 90600 485110
rect 90548 485046 90600 485052
rect 89810 471336 89866 471345
rect 89810 471271 89866 471280
rect 90744 470594 90772 488022
rect 91388 485081 91416 488036
rect 91848 485654 91876 488036
rect 91836 485648 91888 485654
rect 91836 485590 91888 485596
rect 92308 485518 92336 488036
rect 92676 488022 92782 488050
rect 92952 488022 93242 488050
rect 93320 488022 93610 488050
rect 93964 488022 94070 488050
rect 94240 488022 94530 488050
rect 94608 488022 94990 488050
rect 95374 488022 95464 488050
rect 92296 485512 92348 485518
rect 92296 485454 92348 485460
rect 91374 485072 91430 485081
rect 91374 485007 91430 485016
rect 92572 484220 92624 484226
rect 92572 484162 92624 484168
rect 92480 484152 92532 484158
rect 92480 484094 92532 484100
rect 89916 470566 90772 470594
rect 88524 468852 88576 468858
rect 88524 468794 88576 468800
rect 87052 468716 87104 468722
rect 87052 468658 87104 468664
rect 80704 467832 80756 467838
rect 80704 467774 80756 467780
rect 77484 466336 77536 466342
rect 77484 466278 77536 466284
rect 76010 466032 76066 466041
rect 76010 465967 76066 465976
rect 74724 465792 74776 465798
rect 74630 465760 74686 465769
rect 72424 465724 72476 465730
rect 74724 465734 74776 465740
rect 74630 465695 74686 465704
rect 72424 465666 72476 465672
rect 69110 465624 69166 465633
rect 69110 465559 69166 465568
rect 89916 464710 89944 470566
rect 89904 464704 89956 464710
rect 89904 464646 89956 464652
rect 92492 464642 92520 484094
rect 92584 468654 92612 484162
rect 92676 471753 92704 488022
rect 92952 484158 92980 488022
rect 93320 484226 93348 488022
rect 93308 484220 93360 484226
rect 93308 484162 93360 484168
rect 92940 484152 92992 484158
rect 92940 484094 92992 484100
rect 93860 484152 93912 484158
rect 93860 484094 93912 484100
rect 92662 471744 92718 471753
rect 92662 471679 92718 471688
rect 92572 468648 92624 468654
rect 92572 468590 92624 468596
rect 93872 467226 93900 484094
rect 93964 468586 93992 488022
rect 94240 471209 94268 488022
rect 94608 484158 94636 488022
rect 95436 485110 95464 488022
rect 95528 488022 95818 488050
rect 95424 485104 95476 485110
rect 95424 485046 95476 485052
rect 94596 484152 94648 484158
rect 94596 484094 94648 484100
rect 95528 471510 95556 488022
rect 96264 482118 96292 488036
rect 96724 482186 96752 488036
rect 97184 483002 97212 488036
rect 97172 482996 97224 483002
rect 97172 482938 97224 482944
rect 97552 482254 97580 488036
rect 98012 482866 98040 488036
rect 98472 482934 98500 488036
rect 98656 488022 98946 488050
rect 98460 482928 98512 482934
rect 98460 482870 98512 482876
rect 98000 482860 98052 482866
rect 98000 482802 98052 482808
rect 97540 482248 97592 482254
rect 97540 482190 97592 482196
rect 96712 482180 96764 482186
rect 96712 482122 96764 482128
rect 96252 482112 96304 482118
rect 96252 482054 96304 482060
rect 98656 474298 98684 488022
rect 99392 486538 99420 488036
rect 99380 486532 99432 486538
rect 99380 486474 99432 486480
rect 99760 485246 99788 488036
rect 99944 488022 100234 488050
rect 100312 488022 100694 488050
rect 100772 488022 101154 488050
rect 101232 488022 101522 488050
rect 101600 488022 101982 488050
rect 99748 485240 99800 485246
rect 99748 485182 99800 485188
rect 99472 484152 99524 484158
rect 99472 484094 99524 484100
rect 98644 474292 98696 474298
rect 98644 474234 98696 474240
rect 99484 474230 99512 484094
rect 99944 474434 99972 488022
rect 100312 484158 100340 488022
rect 100300 484152 100352 484158
rect 100300 484094 100352 484100
rect 99932 474428 99984 474434
rect 99932 474370 99984 474376
rect 99472 474224 99524 474230
rect 99472 474166 99524 474172
rect 95516 471504 95568 471510
rect 95516 471446 95568 471452
rect 100772 471442 100800 488022
rect 101232 484106 101260 488022
rect 100864 484078 101260 484106
rect 100760 471436 100812 471442
rect 100760 471378 100812 471384
rect 100864 471306 100892 484078
rect 101600 474502 101628 488022
rect 102428 485314 102456 488036
rect 102888 485722 102916 488036
rect 103072 488022 103362 488050
rect 102876 485716 102928 485722
rect 102876 485658 102928 485664
rect 102416 485308 102468 485314
rect 102416 485250 102468 485256
rect 101588 474496 101640 474502
rect 101588 474438 101640 474444
rect 100852 471300 100904 471306
rect 100852 471242 100904 471248
rect 94226 471200 94282 471209
rect 94226 471135 94282 471144
rect 103072 470594 103100 488022
rect 103520 484220 103572 484226
rect 103520 484162 103572 484168
rect 102336 470566 103100 470594
rect 93952 468580 94004 468586
rect 93952 468522 94004 468528
rect 93860 467220 93912 467226
rect 93860 467162 93912 467168
rect 92480 464636 92532 464642
rect 92480 464578 92532 464584
rect 102336 464574 102364 470566
rect 103532 468518 103560 484162
rect 103612 484152 103664 484158
rect 103612 484094 103664 484100
rect 103624 472666 103652 484094
rect 103716 474366 103744 488036
rect 103808 488022 104190 488050
rect 104360 488022 104650 488050
rect 105004 488022 105110 488050
rect 103808 484158 103836 488022
rect 104360 484226 104388 488022
rect 104348 484220 104400 484226
rect 104348 484162 104400 484168
rect 103796 484152 103848 484158
rect 103796 484094 103848 484100
rect 103704 474360 103756 474366
rect 103704 474302 103756 474308
rect 105004 472734 105032 488022
rect 105556 485178 105584 488036
rect 105648 488022 105938 488050
rect 105544 485172 105596 485178
rect 105544 485114 105596 485120
rect 105648 472802 105676 488022
rect 106384 485382 106412 488036
rect 106476 488022 106858 488050
rect 106936 488022 107318 488050
rect 106372 485376 106424 485382
rect 106372 485318 106424 485324
rect 106476 484106 106504 488022
rect 106384 484078 106504 484106
rect 106384 474094 106412 484078
rect 106372 474088 106424 474094
rect 106372 474030 106424 474036
rect 105636 472796 105688 472802
rect 105636 472738 105688 472744
rect 104992 472728 105044 472734
rect 104992 472670 105044 472676
rect 103612 472660 103664 472666
rect 103612 472602 103664 472608
rect 106936 470594 106964 488022
rect 107660 484152 107712 484158
rect 107660 484094 107712 484100
rect 106476 470566 106964 470594
rect 103520 468512 103572 468518
rect 103520 468454 103572 468460
rect 106476 467158 106504 470566
rect 107672 468518 107700 484094
rect 107764 468586 107792 488036
rect 107856 488022 108146 488050
rect 108224 488022 108606 488050
rect 109082 488022 109448 488050
rect 107856 484158 107884 488022
rect 107844 484152 107896 484158
rect 107844 484094 107896 484100
rect 108224 471306 108252 488022
rect 109420 486606 109448 488022
rect 109512 486674 109540 488036
rect 109604 488022 109894 488050
rect 109500 486668 109552 486674
rect 109500 486610 109552 486616
rect 109408 486600 109460 486606
rect 109408 486542 109460 486548
rect 108212 471300 108264 471306
rect 108212 471242 108264 471248
rect 109604 470594 109632 488022
rect 110340 485178 110368 488036
rect 110616 488022 110814 488050
rect 110328 485172 110380 485178
rect 110328 485114 110380 485120
rect 110616 472870 110644 488022
rect 111260 482730 111288 488036
rect 111720 482798 111748 488036
rect 111708 482792 111760 482798
rect 111708 482734 111760 482740
rect 111248 482724 111300 482730
rect 111248 482666 111300 482672
rect 112088 482594 112116 488036
rect 112076 482588 112128 482594
rect 112076 482530 112128 482536
rect 112548 482458 112576 488036
rect 112640 488022 113022 488050
rect 112536 482452 112588 482458
rect 112536 482394 112588 482400
rect 110604 472864 110656 472870
rect 110604 472806 110656 472812
rect 112640 470594 112668 488022
rect 113468 483682 113496 488036
rect 113560 488022 113942 488050
rect 113456 483676 113508 483682
rect 113456 483618 113508 483624
rect 113560 474162 113588 488022
rect 114296 481030 114324 488036
rect 114284 481024 114336 481030
rect 114284 480966 114336 480972
rect 113548 474156 113600 474162
rect 113548 474098 113600 474104
rect 114756 471374 114784 488036
rect 115216 482526 115244 488036
rect 115676 482662 115704 488036
rect 116074 488022 116164 488050
rect 115664 482656 115716 482662
rect 115664 482598 115716 482604
rect 115204 482520 115256 482526
rect 115204 482462 115256 482468
rect 116136 480214 116164 488022
rect 116228 488022 116518 488050
rect 116688 488022 116978 488050
rect 116124 480208 116176 480214
rect 116124 480150 116176 480156
rect 116228 479398 116256 488022
rect 116216 479392 116268 479398
rect 116216 479334 116268 479340
rect 116688 479330 116716 488022
rect 117424 479466 117452 488036
rect 117608 488022 117898 488050
rect 117976 488022 118266 488050
rect 118742 488022 118832 488050
rect 117608 480146 117636 488022
rect 117596 480140 117648 480146
rect 117596 480082 117648 480088
rect 117976 479641 118004 488022
rect 118804 479913 118832 488022
rect 118896 488022 119186 488050
rect 118790 479904 118846 479913
rect 118790 479839 118846 479848
rect 117962 479632 118018 479641
rect 117962 479567 118018 479576
rect 118896 479505 118924 488022
rect 119632 482390 119660 488036
rect 120092 482497 120120 488036
rect 120460 482769 120488 488036
rect 120446 482760 120502 482769
rect 120446 482695 120502 482704
rect 120920 482633 120948 488036
rect 120906 482624 120962 482633
rect 120906 482559 120962 482568
rect 120078 482488 120134 482497
rect 120078 482423 120134 482432
rect 119620 482384 119672 482390
rect 121380 482361 121408 488036
rect 121472 488022 121854 488050
rect 121932 488022 122222 488050
rect 122392 488022 122682 488050
rect 122944 488022 123142 488050
rect 123312 488022 123602 488050
rect 123680 488022 124062 488050
rect 124232 488022 124430 488050
rect 124600 488022 124890 488050
rect 124968 488022 125350 488050
rect 119620 482326 119672 482332
rect 121366 482352 121422 482361
rect 121366 482287 121422 482296
rect 118882 479496 118938 479505
rect 117412 479460 117464 479466
rect 118882 479431 118938 479440
rect 117412 479402 117464 479408
rect 116676 479324 116728 479330
rect 116676 479266 116728 479272
rect 114744 471368 114796 471374
rect 114744 471310 114796 471316
rect 109052 470566 109632 470594
rect 111996 470566 112668 470594
rect 109052 468654 109080 470566
rect 111996 469878 112024 470566
rect 111984 469872 112036 469878
rect 111984 469814 112036 469820
rect 109040 468648 109092 468654
rect 109040 468590 109092 468596
rect 107752 468580 107804 468586
rect 107752 468522 107804 468528
rect 107660 468512 107712 468518
rect 107660 468454 107712 468460
rect 106464 467152 106516 467158
rect 106464 467094 106516 467100
rect 102324 464568 102376 464574
rect 102324 464510 102376 464516
rect 121472 464506 121500 488022
rect 121932 484106 121960 488022
rect 121564 484078 121960 484106
rect 121564 480010 121592 484078
rect 121552 480004 121604 480010
rect 121552 479946 121604 479952
rect 122392 479777 122420 488022
rect 122840 484152 122892 484158
rect 122840 484094 122892 484100
rect 122378 479768 122434 479777
rect 122378 479703 122434 479712
rect 122852 477426 122880 484094
rect 122944 479874 122972 488022
rect 122932 479868 122984 479874
rect 122932 479810 122984 479816
rect 123312 479806 123340 488022
rect 123680 484158 123708 488022
rect 123668 484152 123720 484158
rect 123668 484094 123720 484100
rect 123300 479800 123352 479806
rect 123300 479742 123352 479748
rect 122840 477420 122892 477426
rect 122840 477362 122892 477368
rect 124232 471374 124260 488022
rect 124312 484152 124364 484158
rect 124312 484094 124364 484100
rect 124324 477193 124352 484094
rect 124600 479670 124628 488022
rect 124968 484158 124996 488022
rect 124956 484152 125008 484158
rect 124956 484094 125008 484100
rect 125600 484152 125652 484158
rect 125600 484094 125652 484100
rect 124588 479664 124640 479670
rect 124588 479606 124640 479612
rect 124310 477184 124366 477193
rect 124310 477119 124366 477128
rect 124220 471368 124272 471374
rect 124220 471310 124272 471316
rect 121460 464500 121512 464506
rect 121460 464442 121512 464448
rect 125612 464409 125640 484094
rect 125692 482044 125744 482050
rect 125692 481986 125744 481992
rect 125704 477057 125732 481986
rect 125690 477048 125746 477057
rect 125690 476983 125746 476992
rect 125796 476921 125824 488036
rect 125888 488022 126270 488050
rect 126348 488022 126638 488050
rect 126992 488022 127098 488050
rect 127176 488022 127558 488050
rect 127728 488022 128018 488050
rect 128372 488022 128478 488050
rect 128556 488022 128846 488050
rect 129016 488022 129306 488050
rect 125888 482050 125916 488022
rect 126348 484158 126376 488022
rect 126336 484152 126388 484158
rect 126336 484094 126388 484100
rect 125876 482044 125928 482050
rect 125876 481986 125928 481992
rect 125782 476912 125838 476921
rect 125782 476847 125838 476856
rect 126992 464506 127020 488022
rect 127176 484106 127204 488022
rect 127084 484078 127204 484106
rect 127084 476785 127112 484078
rect 127728 479942 127756 488022
rect 127716 479936 127768 479942
rect 127716 479878 127768 479884
rect 127070 476776 127126 476785
rect 127070 476711 127126 476720
rect 126980 464500 127032 464506
rect 126980 464442 127032 464448
rect 128372 464438 128400 488022
rect 128556 484106 128584 488022
rect 128464 484078 128584 484106
rect 128464 476610 128492 484078
rect 129016 479602 129044 488022
rect 129752 479738 129780 488036
rect 130028 488022 130226 488050
rect 130304 488022 130594 488050
rect 130672 488022 131054 488050
rect 131316 488022 131514 488050
rect 131592 488022 131974 488050
rect 132144 488022 132434 488050
rect 132512 488022 132802 488050
rect 132880 488022 133262 488050
rect 133432 488022 133722 488050
rect 133984 488022 134182 488050
rect 134352 488022 134642 488050
rect 134720 488022 135010 488050
rect 135486 488022 135760 488050
rect 129832 484220 129884 484226
rect 129832 484162 129884 484168
rect 129740 479732 129792 479738
rect 129740 479674 129792 479680
rect 129004 479596 129056 479602
rect 129004 479538 129056 479544
rect 129844 477154 129872 484162
rect 129924 484152 129976 484158
rect 129924 484094 129976 484100
rect 129936 480078 129964 484094
rect 129924 480072 129976 480078
rect 129924 480014 129976 480020
rect 129832 477148 129884 477154
rect 129832 477090 129884 477096
rect 128452 476604 128504 476610
rect 128452 476546 128504 476552
rect 128360 464432 128412 464438
rect 125598 464400 125654 464409
rect 128360 464374 128412 464380
rect 130028 464370 130056 488022
rect 130304 484158 130332 488022
rect 130672 484226 130700 488022
rect 130660 484220 130712 484226
rect 130660 484162 130712 484168
rect 130292 484152 130344 484158
rect 130292 484094 130344 484100
rect 131120 484152 131172 484158
rect 131120 484094 131172 484100
rect 131132 476678 131160 484094
rect 131212 480684 131264 480690
rect 131212 480626 131264 480632
rect 131224 476746 131252 480626
rect 131316 477222 131344 488022
rect 131592 480690 131620 488022
rect 132144 484158 132172 488022
rect 132132 484152 132184 484158
rect 132132 484094 132184 484100
rect 131580 480684 131632 480690
rect 131580 480626 131632 480632
rect 131304 477216 131356 477222
rect 131304 477158 131356 477164
rect 132512 476950 132540 488022
rect 132880 484106 132908 488022
rect 132604 484078 132908 484106
rect 132604 477018 132632 484078
rect 133432 477086 133460 488022
rect 133880 484152 133932 484158
rect 133880 484094 133932 484100
rect 133892 477494 133920 484094
rect 133880 477488 133932 477494
rect 133880 477430 133932 477436
rect 133420 477080 133472 477086
rect 133420 477022 133472 477028
rect 132592 477012 132644 477018
rect 132592 476954 132644 476960
rect 132500 476944 132552 476950
rect 132500 476886 132552 476892
rect 133984 476882 134012 488022
rect 134352 484158 134380 488022
rect 134340 484152 134392 484158
rect 134340 484094 134392 484100
rect 134720 477290 134748 488022
rect 135732 482526 135760 488022
rect 135720 482520 135772 482526
rect 135720 482462 135772 482468
rect 135916 482322 135944 488036
rect 136008 488022 136390 488050
rect 136652 488022 136758 488050
rect 137234 488022 137600 488050
rect 137694 488022 137968 488050
rect 138154 488022 138520 488050
rect 138614 488022 138888 488050
rect 138982 488022 139256 488050
rect 135904 482316 135956 482322
rect 135904 482258 135956 482264
rect 136008 477358 136036 488022
rect 135996 477352 136048 477358
rect 135996 477294 136048 477300
rect 134708 477284 134760 477290
rect 134708 477226 134760 477232
rect 133972 476876 134024 476882
rect 133972 476818 134024 476824
rect 131212 476740 131264 476746
rect 131212 476682 131264 476688
rect 131120 476672 131172 476678
rect 131120 476614 131172 476620
rect 136652 464370 136680 488022
rect 137572 482322 137600 488022
rect 137940 482390 137968 488022
rect 138492 482662 138520 488022
rect 138480 482656 138532 482662
rect 138480 482598 138532 482604
rect 138860 482458 138888 488022
rect 139228 485246 139256 488022
rect 139216 485240 139268 485246
rect 139216 485182 139268 485188
rect 139412 484906 139440 488036
rect 139504 488022 139886 488050
rect 140056 488022 140346 488050
rect 140822 488022 140912 488050
rect 139400 484900 139452 484906
rect 139400 484842 139452 484848
rect 139400 484152 139452 484158
rect 139400 484094 139452 484100
rect 138848 482452 138900 482458
rect 138848 482394 138900 482400
rect 137928 482384 137980 482390
rect 137928 482326 137980 482332
rect 137560 482316 137612 482322
rect 137560 482258 137612 482264
rect 139412 468722 139440 484094
rect 139504 474094 139532 488022
rect 140056 484158 140084 488022
rect 140884 486538 140912 488022
rect 140976 488022 141174 488050
rect 141344 488022 141634 488050
rect 141712 488022 142094 488050
rect 142264 488022 142554 488050
rect 142632 488022 142922 488050
rect 143000 488022 143382 488050
rect 140872 486532 140924 486538
rect 140872 486474 140924 486480
rect 140044 484152 140096 484158
rect 140044 484094 140096 484100
rect 140872 484152 140924 484158
rect 140872 484094 140924 484100
rect 140780 482588 140832 482594
rect 140780 482530 140832 482536
rect 139492 474088 139544 474094
rect 139492 474030 139544 474036
rect 139400 468716 139452 468722
rect 139400 468658 139452 468664
rect 140792 465866 140820 482530
rect 140884 471442 140912 484094
rect 140976 471510 141004 488022
rect 141344 482594 141372 488022
rect 141712 484158 141740 488022
rect 141700 484152 141752 484158
rect 141700 484094 141752 484100
rect 142160 484152 142212 484158
rect 142160 484094 142212 484100
rect 141332 482588 141384 482594
rect 141332 482530 141384 482536
rect 140964 471504 141016 471510
rect 140964 471446 141016 471452
rect 140872 471436 140924 471442
rect 140872 471378 140924 471384
rect 140780 465860 140832 465866
rect 140780 465802 140832 465808
rect 142172 464438 142200 484094
rect 142264 465798 142292 488022
rect 142632 484158 142660 488022
rect 142620 484152 142672 484158
rect 142620 484094 142672 484100
rect 143000 470594 143028 488022
rect 143632 484220 143684 484226
rect 143632 484162 143684 484168
rect 143540 484152 143592 484158
rect 143540 484094 143592 484100
rect 143552 472569 143580 484094
rect 143644 474065 143672 484162
rect 143828 480298 143856 488036
rect 143920 488022 144302 488050
rect 144472 488022 144762 488050
rect 145146 488022 145512 488050
rect 145606 488022 145696 488050
rect 143920 484226 143948 488022
rect 143908 484220 143960 484226
rect 143908 484162 143960 484168
rect 144472 484158 144500 488022
rect 145484 485081 145512 488022
rect 145668 485353 145696 488022
rect 145760 488022 146050 488050
rect 146312 488022 146510 488050
rect 146986 488022 147260 488050
rect 147354 488022 147628 488050
rect 145654 485344 145710 485353
rect 145654 485279 145710 485288
rect 145470 485072 145526 485081
rect 145470 485007 145526 485016
rect 144460 484152 144512 484158
rect 144460 484094 144512 484100
rect 143736 480270 143856 480298
rect 143736 476814 143764 480270
rect 145760 476921 145788 488022
rect 146312 478174 146340 488022
rect 147232 480865 147260 488022
rect 147600 485217 147628 488022
rect 147586 485208 147642 485217
rect 147586 485143 147642 485152
rect 147680 484152 147732 484158
rect 147680 484094 147732 484100
rect 147218 480856 147274 480865
rect 147218 480791 147274 480800
rect 146300 478168 146352 478174
rect 146300 478110 146352 478116
rect 145746 476912 145802 476921
rect 145746 476847 145802 476856
rect 143724 476808 143776 476814
rect 143724 476750 143776 476756
rect 143630 474056 143686 474065
rect 143630 473991 143686 474000
rect 143538 472560 143594 472569
rect 143538 472495 143594 472504
rect 142356 470566 143028 470594
rect 142356 468790 142384 470566
rect 147692 469849 147720 484094
rect 147784 479641 147812 488036
rect 148244 485314 148272 488036
rect 148336 488022 148718 488050
rect 149194 488022 149468 488050
rect 149562 488022 149928 488050
rect 150022 488022 150296 488050
rect 148232 485308 148284 485314
rect 148232 485250 148284 485256
rect 148336 484158 148364 488022
rect 149440 485450 149468 488022
rect 149428 485444 149480 485450
rect 149428 485386 149480 485392
rect 149900 485042 149928 488022
rect 149888 485036 149940 485042
rect 149888 484978 149940 484984
rect 148324 484152 148376 484158
rect 148324 484094 148376 484100
rect 150268 483721 150296 488022
rect 150452 485586 150480 488036
rect 150544 488022 150926 488050
rect 150440 485580 150492 485586
rect 150440 485522 150492 485528
rect 150544 484140 150572 488022
rect 151280 485790 151308 488036
rect 151372 488022 151754 488050
rect 151268 485784 151320 485790
rect 151268 485726 151320 485732
rect 150452 484112 150572 484140
rect 150254 483712 150310 483721
rect 150254 483647 150310 483656
rect 147770 479632 147826 479641
rect 147770 479567 147826 479576
rect 150452 475425 150480 484112
rect 151372 476785 151400 488022
rect 152200 485518 152228 488036
rect 152292 488022 152674 488050
rect 152752 488022 153134 488050
rect 153212 488022 153502 488050
rect 152188 485512 152240 485518
rect 152188 485454 152240 485460
rect 152292 484106 152320 488022
rect 151832 484078 152320 484106
rect 151358 476776 151414 476785
rect 151358 476711 151414 476720
rect 150438 475416 150494 475425
rect 150438 475351 150494 475360
rect 147678 469840 147734 469849
rect 147678 469775 147734 469784
rect 142344 468784 142396 468790
rect 142344 468726 142396 468732
rect 151832 467158 151860 484078
rect 152752 478281 152780 488022
rect 152738 478272 152794 478281
rect 152738 478207 152794 478216
rect 153212 474162 153240 488022
rect 153948 485722 153976 488036
rect 154040 488022 154422 488050
rect 154898 488022 155264 488050
rect 155358 488022 155632 488050
rect 155726 488022 155908 488050
rect 156186 488022 156552 488050
rect 153936 485716 153988 485722
rect 153936 485658 153988 485664
rect 154040 479505 154068 488022
rect 155236 481001 155264 488022
rect 155604 484770 155632 488022
rect 155592 484764 155644 484770
rect 155592 484706 155644 484712
rect 155880 482361 155908 488022
rect 156524 483857 156552 488022
rect 156616 484974 156644 488036
rect 156708 488022 157090 488050
rect 156604 484968 156656 484974
rect 156604 484910 156656 484916
rect 156510 483848 156566 483857
rect 156510 483783 156566 483792
rect 155866 482352 155922 482361
rect 155866 482287 155922 482296
rect 155222 480992 155278 481001
rect 155222 480927 155278 480936
rect 154026 479496 154082 479505
rect 154026 479431 154082 479440
rect 153200 474156 153252 474162
rect 153200 474098 153252 474104
rect 156708 470594 156736 488022
rect 157444 484838 157472 488036
rect 157536 488022 157918 488050
rect 158394 488022 158668 488050
rect 157432 484832 157484 484838
rect 157432 484774 157484 484780
rect 157536 475561 157564 488022
rect 158640 485761 158668 488022
rect 158732 488022 158838 488050
rect 159008 488022 159298 488050
rect 159682 488022 160048 488050
rect 160142 488022 160232 488050
rect 158626 485752 158682 485761
rect 158626 485687 158682 485696
rect 157522 475552 157578 475561
rect 157522 475487 157578 475496
rect 158732 474230 158760 488022
rect 159008 479602 159036 488022
rect 160020 483682 160048 488022
rect 160100 484152 160152 484158
rect 160100 484094 160152 484100
rect 160008 483676 160060 483682
rect 160008 483618 160060 483624
rect 158996 479596 159048 479602
rect 158996 479538 159048 479544
rect 158720 474224 158772 474230
rect 158720 474166 158772 474172
rect 155972 470566 156736 470594
rect 151820 467152 151872 467158
rect 155972 467129 156000 470566
rect 160112 469878 160140 484094
rect 160204 478242 160232 488022
rect 160572 481030 160600 488036
rect 160664 488022 161046 488050
rect 161522 488022 161612 488050
rect 160664 484158 160692 488022
rect 161584 484294 161612 488022
rect 161676 488022 161874 488050
rect 161952 488022 162334 488050
rect 162504 488022 162794 488050
rect 162964 488022 163254 488050
rect 163638 488022 163728 488050
rect 161572 484288 161624 484294
rect 161572 484230 161624 484236
rect 161480 484220 161532 484226
rect 161480 484162 161532 484168
rect 160652 484152 160704 484158
rect 160652 484094 160704 484100
rect 160560 481024 160612 481030
rect 160560 480966 160612 480972
rect 160192 478236 160244 478242
rect 160192 478178 160244 478184
rect 160100 469872 160152 469878
rect 160100 469814 160152 469820
rect 161492 468489 161520 484162
rect 161572 484152 161624 484158
rect 161572 484094 161624 484100
rect 161584 471345 161612 484094
rect 161676 471578 161704 488022
rect 161952 484226 161980 488022
rect 161940 484220 161992 484226
rect 161940 484162 161992 484168
rect 162504 484158 162532 488022
rect 162768 484288 162820 484294
rect 162768 484230 162820 484236
rect 162492 484152 162544 484158
rect 162492 484094 162544 484100
rect 162780 483750 162808 484230
rect 162860 484152 162912 484158
rect 162860 484094 162912 484100
rect 162768 483744 162820 483750
rect 162768 483686 162820 483692
rect 161664 471572 161716 471578
rect 161664 471514 161716 471520
rect 161570 471336 161626 471345
rect 161570 471271 161626 471280
rect 161478 468480 161534 468489
rect 161478 468415 161534 468424
rect 151820 467094 151872 467100
rect 155958 467120 156014 467129
rect 155958 467055 156014 467064
rect 162872 465905 162900 484094
rect 162964 475522 162992 488022
rect 163700 485489 163728 488022
rect 163792 488022 164082 488050
rect 164252 488022 164542 488050
rect 164620 488022 165002 488050
rect 165478 488022 165568 488050
rect 163686 485480 163742 485489
rect 163686 485415 163742 485424
rect 163792 484158 163820 488022
rect 163780 484152 163832 484158
rect 163780 484094 163832 484100
rect 162952 475516 163004 475522
rect 162952 475458 163004 475464
rect 164252 467226 164280 488022
rect 164620 476814 164648 488022
rect 164884 485172 164936 485178
rect 164884 485114 164936 485120
rect 164608 476808 164660 476814
rect 164608 476750 164660 476756
rect 164240 467220 164292 467226
rect 164240 467162 164292 467168
rect 164896 466002 164924 485114
rect 165540 482662 165568 488022
rect 165632 488022 165830 488050
rect 165528 482656 165580 482662
rect 165528 482598 165580 482604
rect 164884 465996 164936 466002
rect 164884 465938 164936 465944
rect 162858 465896 162914 465905
rect 162858 465831 162914 465840
rect 142252 465792 142304 465798
rect 165632 465769 165660 488022
rect 166172 485648 166224 485654
rect 166172 485590 166224 485596
rect 166184 484974 166212 485590
rect 166276 485178 166304 488036
rect 166368 488022 166750 488050
rect 167012 488022 167210 488050
rect 167288 488022 167670 488050
rect 167748 488022 168038 488050
rect 168514 488022 168604 488050
rect 166264 485172 166316 485178
rect 166264 485114 166316 485120
rect 166172 484968 166224 484974
rect 166172 484910 166224 484916
rect 166264 484968 166316 484974
rect 166264 484910 166316 484916
rect 166276 484770 166304 484910
rect 166264 484764 166316 484770
rect 166264 484706 166316 484712
rect 166368 470594 166396 488022
rect 165816 470566 166396 470594
rect 165816 466177 165844 470566
rect 165802 466168 165858 466177
rect 165802 466103 165858 466112
rect 167012 466041 167040 488022
rect 167092 480888 167144 480894
rect 167092 480830 167144 480836
rect 167104 468897 167132 480830
rect 167288 470594 167316 488022
rect 167748 480894 167776 488022
rect 167828 485104 167880 485110
rect 167828 485046 167880 485052
rect 167840 484770 167868 485046
rect 167828 484764 167880 484770
rect 167828 484706 167880 484712
rect 168576 481098 168604 488022
rect 168668 488022 168958 488050
rect 169128 488022 169418 488050
rect 169894 488022 169984 488050
rect 168564 481092 168616 481098
rect 168564 481034 168616 481040
rect 167736 480888 167788 480894
rect 167736 480830 167788 480836
rect 168380 480888 168432 480894
rect 168380 480830 168432 480836
rect 167196 470566 167316 470594
rect 167090 468888 167146 468897
rect 167196 468858 167224 470566
rect 167090 468823 167146 468832
rect 167184 468852 167236 468858
rect 167184 468794 167236 468800
rect 168392 468625 168420 480830
rect 168668 475454 168696 488022
rect 168748 481092 168800 481098
rect 168748 481034 168800 481040
rect 168656 475448 168708 475454
rect 168656 475390 168708 475396
rect 168760 473354 168788 481034
rect 169128 480894 169156 488022
rect 169116 480888 169168 480894
rect 169116 480830 169168 480836
rect 169760 480888 169812 480894
rect 169760 480830 169812 480836
rect 168576 473326 168788 473354
rect 168576 468761 168604 473326
rect 169772 471617 169800 480830
rect 169852 478780 169904 478786
rect 169852 478722 169904 478728
rect 169864 472705 169892 478722
rect 169850 472696 169906 472705
rect 169850 472631 169906 472640
rect 169956 471753 169984 488022
rect 170048 488022 170246 488050
rect 170416 488022 170706 488050
rect 170048 480894 170076 488022
rect 170036 480888 170088 480894
rect 170036 480830 170088 480836
rect 170416 478786 170444 488022
rect 171152 485625 171180 488036
rect 171244 488022 171626 488050
rect 171704 488022 171994 488050
rect 172072 488022 172454 488050
rect 172532 488022 172914 488050
rect 173390 488022 173480 488050
rect 171138 485616 171194 485625
rect 171138 485551 171194 485560
rect 171140 480344 171192 480350
rect 171140 480286 171192 480292
rect 170404 478780 170456 478786
rect 170404 478722 170456 478728
rect 169942 471744 169998 471753
rect 169942 471679 169998 471688
rect 169758 471608 169814 471617
rect 169758 471543 169814 471552
rect 171152 471209 171180 480286
rect 171244 472841 171272 488022
rect 171704 480350 171732 488022
rect 171692 480344 171744 480350
rect 171692 480286 171744 480292
rect 172072 474298 172100 488022
rect 172060 474292 172112 474298
rect 172060 474234 172112 474240
rect 171230 472832 171286 472841
rect 171230 472767 171286 472776
rect 171138 471200 171194 471209
rect 171138 471135 171194 471144
rect 172532 469033 172560 488022
rect 173452 482730 173480 488022
rect 173544 488022 173834 488050
rect 174004 488022 174202 488050
rect 174280 488022 174662 488050
rect 174832 488022 175122 488050
rect 175384 488022 175582 488050
rect 173440 482724 173492 482730
rect 173440 482666 173492 482672
rect 173544 470594 173572 488022
rect 173900 480888 173952 480894
rect 173900 480830 173952 480836
rect 172624 470566 173572 470594
rect 172624 469946 172652 470566
rect 172612 469940 172664 469946
rect 172612 469882 172664 469888
rect 172518 469024 172574 469033
rect 172518 468959 172574 468968
rect 168562 468752 168618 468761
rect 168562 468687 168618 468696
rect 168378 468616 168434 468625
rect 168378 468551 168434 468560
rect 166998 466032 167054 466041
rect 166998 465967 167054 465976
rect 173912 465934 173940 480830
rect 174004 466138 174032 488022
rect 174280 480894 174308 488022
rect 174268 480888 174320 480894
rect 174268 480830 174320 480836
rect 174832 471481 174860 488022
rect 175280 476468 175332 476474
rect 175280 476410 175332 476416
rect 174818 471472 174874 471481
rect 174818 471407 174874 471416
rect 175292 469062 175320 476410
rect 175384 472734 175412 488022
rect 176028 481098 176056 488036
rect 176120 488022 176410 488050
rect 176886 488022 177160 488050
rect 176016 481092 176068 481098
rect 176016 481034 176068 481040
rect 176120 476474 176148 488022
rect 177132 482798 177160 488022
rect 177316 483818 177344 488036
rect 177408 488022 177790 488050
rect 177304 483812 177356 483818
rect 177304 483754 177356 483760
rect 177120 482792 177172 482798
rect 177120 482734 177172 482740
rect 176108 476468 176160 476474
rect 176108 476410 176160 476416
rect 175372 472728 175424 472734
rect 175372 472670 175424 472676
rect 177408 470594 177436 488022
rect 178144 478310 178172 488036
rect 178328 488022 178618 488050
rect 178696 488022 179078 488050
rect 178132 478304 178184 478310
rect 178132 478246 178184 478252
rect 178328 476114 178356 488022
rect 178696 479777 178724 488022
rect 179420 480888 179472 480894
rect 179420 480830 179472 480836
rect 178682 479768 178738 479777
rect 178682 479703 178738 479712
rect 178052 476086 178356 476114
rect 178052 474366 178080 476086
rect 178040 474360 178092 474366
rect 178040 474302 178092 474308
rect 176672 470566 177436 470594
rect 175280 469056 175332 469062
rect 175280 468998 175332 469004
rect 173992 466132 174044 466138
rect 173992 466074 174044 466080
rect 176672 466070 176700 470566
rect 179432 468926 179460 480830
rect 179524 472666 179552 488036
rect 179616 488022 179998 488050
rect 180076 488022 180366 488050
rect 179616 475590 179644 488022
rect 180076 480894 180104 488022
rect 180064 480888 180116 480894
rect 180064 480830 180116 480836
rect 179604 475584 179656 475590
rect 179604 475526 179656 475532
rect 180156 474020 180208 474026
rect 180156 473962 180208 473968
rect 179512 472660 179564 472666
rect 179512 472602 179564 472608
rect 179420 468920 179472 468926
rect 179420 468862 179472 468868
rect 178040 467832 178092 467838
rect 178040 467774 178092 467780
rect 178052 466585 178080 467774
rect 180168 467294 180196 473962
rect 180156 467288 180208 467294
rect 180154 467256 180156 467265
rect 180208 467256 180210 467265
rect 180154 467191 180210 467200
rect 178038 466576 178094 466585
rect 178038 466511 178040 466520
rect 178092 466511 178094 466520
rect 178040 466482 178092 466488
rect 178052 466451 178080 466482
rect 180812 466206 180840 488036
rect 180904 488022 181286 488050
rect 181456 488022 181746 488050
rect 180904 468994 180932 488022
rect 181456 471782 181484 488022
rect 181444 471776 181496 471782
rect 181444 471718 181496 471724
rect 180892 468988 180944 468994
rect 180892 468930 180944 468936
rect 182192 466410 182220 488036
rect 182376 488022 182574 488050
rect 182744 488022 183034 488050
rect 183112 488022 183494 488050
rect 183572 488022 183954 488050
rect 184032 488022 184322 488050
rect 184798 488022 184888 488050
rect 182270 485752 182326 485761
rect 182270 485687 182326 485696
rect 182284 485110 182312 485687
rect 182272 485104 182324 485110
rect 182272 485046 182324 485052
rect 182272 480888 182324 480894
rect 182272 480830 182324 480836
rect 182284 471646 182312 480830
rect 182272 471640 182324 471646
rect 182272 471582 182324 471588
rect 182376 471238 182404 488022
rect 182744 471714 182772 488022
rect 182824 484764 182876 484770
rect 182824 484706 182876 484712
rect 182732 471708 182784 471714
rect 182732 471650 182784 471656
rect 182364 471232 182416 471238
rect 182364 471174 182416 471180
rect 182180 466404 182232 466410
rect 182180 466346 182232 466352
rect 182836 466313 182864 484706
rect 183112 480894 183140 488022
rect 183100 480888 183152 480894
rect 183100 480830 183152 480836
rect 182822 466304 182878 466313
rect 182822 466239 182878 466248
rect 180800 466200 180852 466206
rect 180800 466142 180852 466148
rect 176660 466064 176712 466070
rect 176660 466006 176712 466012
rect 173900 465928 173952 465934
rect 173900 465870 173952 465876
rect 142252 465734 142304 465740
rect 165618 465760 165674 465769
rect 165618 465695 165674 465704
rect 183572 464642 183600 488022
rect 184032 470594 184060 488022
rect 184860 485761 184888 488022
rect 184952 488022 185242 488050
rect 185320 488022 185702 488050
rect 185780 488022 186162 488050
rect 186424 488022 186530 488050
rect 187006 488022 187096 488050
rect 184846 485752 184902 485761
rect 184846 485687 184902 485696
rect 183664 470566 184060 470594
rect 183664 464710 183692 470566
rect 184952 467362 184980 488022
rect 185320 476114 185348 488022
rect 185584 484900 185636 484906
rect 185584 484842 185636 484848
rect 185044 476086 185348 476114
rect 185044 471986 185072 476086
rect 185032 471980 185084 471986
rect 185032 471922 185084 471928
rect 185596 471170 185624 484842
rect 185780 476882 185808 488022
rect 186320 485376 186372 485382
rect 186320 485318 186372 485324
rect 186332 485246 186360 485318
rect 186320 485240 186372 485246
rect 186320 485182 186372 485188
rect 186320 480888 186372 480894
rect 186320 480830 186372 480836
rect 185768 476876 185820 476882
rect 185768 476818 185820 476824
rect 185584 471164 185636 471170
rect 185584 471106 185636 471112
rect 186332 468314 186360 480830
rect 186424 474026 186452 488022
rect 187068 484945 187096 488022
rect 187160 488022 187450 488050
rect 187712 488022 187910 488050
rect 188080 488022 188370 488050
rect 188448 488022 188738 488050
rect 187054 484936 187110 484945
rect 187054 484871 187110 484880
rect 187160 480894 187188 488022
rect 187148 480888 187200 480894
rect 187148 480830 187200 480836
rect 186412 474020 186464 474026
rect 186412 473962 186464 473968
rect 186320 468308 186372 468314
rect 186320 468250 186372 468256
rect 184940 467356 184992 467362
rect 184940 467298 184992 467304
rect 187712 466342 187740 488022
rect 188080 476950 188108 488022
rect 188068 476944 188120 476950
rect 188068 476886 188120 476892
rect 188448 476114 188476 488022
rect 189184 481166 189212 488036
rect 189368 488022 189658 488050
rect 189736 488022 190118 488050
rect 189368 485774 189396 488022
rect 189276 485746 189396 485774
rect 189172 481160 189224 481166
rect 189172 481102 189224 481108
rect 189276 478122 189304 485746
rect 189356 481160 189408 481166
rect 189356 481102 189408 481108
rect 187804 476086 188476 476114
rect 189092 478094 189304 478122
rect 187804 475658 187832 476086
rect 187792 475652 187844 475658
rect 187792 475594 187844 475600
rect 189092 467430 189120 478094
rect 189368 473354 189396 481102
rect 189184 473326 189396 473354
rect 189184 467498 189212 473326
rect 189736 471918 189764 488022
rect 189724 471912 189776 471918
rect 189724 471854 189776 471860
rect 189172 467492 189224 467498
rect 189172 467434 189224 467440
rect 189080 467424 189132 467430
rect 189080 467366 189132 467372
rect 187700 466336 187752 466342
rect 187700 466278 187752 466284
rect 190472 464778 190500 488036
rect 190564 488022 190946 488050
rect 191024 488022 191406 488050
rect 190564 465662 190592 488022
rect 191024 471850 191052 488022
rect 191196 485444 191248 485450
rect 191196 485386 191248 485392
rect 191102 485208 191158 485217
rect 191102 485143 191158 485152
rect 191116 484673 191144 485143
rect 191208 484906 191236 485386
rect 191196 484900 191248 484906
rect 191196 484842 191248 484848
rect 191102 484664 191158 484673
rect 191102 484599 191158 484608
rect 191012 471844 191064 471850
rect 191012 471786 191064 471792
rect 190918 466576 190974 466585
rect 190918 466511 190974 466520
rect 190932 466478 190960 466511
rect 190920 466472 190972 466478
rect 190920 466414 190972 466420
rect 191852 466274 191880 488036
rect 191944 488022 192326 488050
rect 192404 488022 192694 488050
rect 192864 488022 193154 488050
rect 193232 488022 193614 488050
rect 193692 488022 194074 488050
rect 194152 488022 194534 488050
rect 194918 488022 195192 488050
rect 191944 468450 191972 488022
rect 192404 476114 192432 488022
rect 192036 476086 192432 476114
rect 192036 469198 192064 476086
rect 192864 470594 192892 488022
rect 192128 470566 192892 470594
rect 192024 469192 192076 469198
rect 192024 469134 192076 469140
rect 191932 468444 191984 468450
rect 191932 468386 191984 468392
rect 192128 468382 192156 470566
rect 192116 468376 192168 468382
rect 192116 468318 192168 468324
rect 191840 466268 191892 466274
rect 191840 466210 191892 466216
rect 190552 465656 190604 465662
rect 190552 465598 190604 465604
rect 190460 464772 190512 464778
rect 190460 464714 190512 464720
rect 183652 464704 183704 464710
rect 183652 464646 183704 464652
rect 183560 464636 183612 464642
rect 183560 464578 183612 464584
rect 193232 464574 193260 488022
rect 193692 476114 193720 488022
rect 194152 485774 194180 488022
rect 193324 476086 193720 476114
rect 193784 485746 194180 485774
rect 193324 465526 193352 476086
rect 193784 470594 193812 485746
rect 193864 485376 193916 485382
rect 193864 485318 193916 485324
rect 193876 471034 193904 485318
rect 195164 484430 195192 488022
rect 195256 488022 195362 488050
rect 195440 488022 195822 488050
rect 196298 488022 196664 488050
rect 196758 488022 196848 488050
rect 195256 485314 195284 488022
rect 195244 485308 195296 485314
rect 195244 485250 195296 485256
rect 195152 484424 195204 484430
rect 195152 484366 195204 484372
rect 195244 471436 195296 471442
rect 195244 471378 195296 471384
rect 195336 471436 195388 471442
rect 195336 471378 195388 471384
rect 195256 471102 195284 471378
rect 195244 471096 195296 471102
rect 195244 471038 195296 471044
rect 195348 471034 195376 471378
rect 193864 471028 193916 471034
rect 193864 470970 193916 470976
rect 195336 471028 195388 471034
rect 195336 470970 195388 470976
rect 195440 470594 195468 488022
rect 193416 470566 193812 470594
rect 194612 470566 195468 470594
rect 193416 469130 193444 470566
rect 193404 469124 193456 469130
rect 193404 469066 193456 469072
rect 194612 465594 194640 470566
rect 194600 465588 194652 465594
rect 194600 465530 194652 465536
rect 193312 465520 193364 465526
rect 193312 465462 193364 465468
rect 193220 464568 193272 464574
rect 193220 464510 193272 464516
rect 142160 464432 142212 464438
rect 142160 464374 142212 464380
rect 125598 464335 125654 464344
rect 130016 464364 130068 464370
rect 130016 464306 130068 464312
rect 136640 464364 136692 464370
rect 136640 464306 136692 464312
rect 196532 381064 196584 381070
rect 60002 381032 60058 381041
rect 196532 381006 196584 381012
rect 60002 380967 60058 380976
rect 59912 166524 59964 166530
rect 59912 166466 59964 166472
rect 59820 165572 59872 165578
rect 59820 165514 59872 165520
rect 59912 164212 59964 164218
rect 59912 164154 59964 164160
rect 59452 164008 59504 164014
rect 59452 163950 59504 163956
rect 59464 163538 59492 163950
rect 59924 163674 59952 164154
rect 59912 163668 59964 163674
rect 59912 163610 59964 163616
rect 59452 163532 59504 163538
rect 59452 163474 59504 163480
rect 59360 146260 59412 146266
rect 59360 146202 59412 146208
rect 59372 146062 59400 146202
rect 59360 146056 59412 146062
rect 59360 145998 59412 146004
rect 59464 140865 59492 163474
rect 59820 148572 59872 148578
rect 59820 148514 59872 148520
rect 59728 146124 59780 146130
rect 59728 146066 59780 146072
rect 59450 140856 59506 140865
rect 59450 140791 59506 140800
rect 59740 59294 59768 146066
rect 59728 59288 59780 59294
rect 59728 59230 59780 59236
rect 59832 58886 59860 148514
rect 59820 58880 59872 58886
rect 59820 58822 59872 58828
rect 59268 57316 59320 57322
rect 59268 57258 59320 57264
rect 59924 55010 59952 163610
rect 60016 57458 60044 380967
rect 60096 380928 60148 380934
rect 143540 380928 143592 380934
rect 60096 380870 60148 380876
rect 93398 380896 93454 380905
rect 60108 358086 60136 380870
rect 93398 380831 93454 380840
rect 110970 380896 111026 380905
rect 110970 380831 111026 380840
rect 113546 380896 113602 380905
rect 113546 380831 113602 380840
rect 116030 380896 116086 380905
rect 116030 380831 116086 380840
rect 118422 380896 118478 380905
rect 118422 380831 118478 380840
rect 120998 380896 121054 380905
rect 120998 380831 121054 380840
rect 123482 380896 123538 380905
rect 123482 380831 123538 380840
rect 125966 380896 126022 380905
rect 125966 380831 126022 380840
rect 131026 380896 131082 380905
rect 131026 380831 131082 380840
rect 133510 380896 133566 380905
rect 133510 380831 133566 380840
rect 135902 380896 135958 380905
rect 135902 380831 135958 380840
rect 143538 380896 143540 380905
rect 143592 380896 143594 380905
rect 143538 380831 143594 380840
rect 146022 380896 146078 380905
rect 146022 380831 146078 380840
rect 158534 380896 158590 380905
rect 158534 380831 158590 380840
rect 160926 380896 160982 380905
rect 160926 380831 160982 380840
rect 163410 380896 163466 380905
rect 163410 380831 163466 380840
rect 165986 380896 166042 380905
rect 165986 380831 166042 380840
rect 87696 379500 87748 379506
rect 87696 379442 87748 379448
rect 87708 379409 87736 379442
rect 85486 379400 85542 379409
rect 85486 379335 85542 379344
rect 86590 379400 86646 379409
rect 86590 379335 86646 379344
rect 87694 379400 87750 379409
rect 87694 379335 87750 379344
rect 88338 379400 88394 379409
rect 88338 379335 88340 379344
rect 80426 379264 80482 379273
rect 80426 379199 80482 379208
rect 81438 379264 81494 379273
rect 81438 379199 81494 379208
rect 80440 378457 80468 379199
rect 80426 378448 80482 378457
rect 80426 378383 80482 378392
rect 80440 378214 80468 378383
rect 81452 378282 81480 379199
rect 83462 378856 83518 378865
rect 83462 378791 83518 378800
rect 81440 378276 81492 378282
rect 81440 378218 81492 378224
rect 80428 378208 80480 378214
rect 80428 378150 80480 378156
rect 83476 376650 83504 378791
rect 85500 378214 85528 379335
rect 86604 378690 86632 379335
rect 88392 379335 88394 379344
rect 88798 379400 88854 379409
rect 88798 379335 88800 379344
rect 88340 379306 88392 379312
rect 88852 379335 88854 379344
rect 90086 379400 90142 379409
rect 90086 379335 90142 379344
rect 90638 379400 90694 379409
rect 90638 379335 90694 379344
rect 91374 379400 91430 379409
rect 91374 379335 91430 379344
rect 92386 379400 92442 379409
rect 92386 379335 92442 379344
rect 88800 379306 88852 379312
rect 90100 378826 90128 379335
rect 90652 379302 90680 379335
rect 91388 379302 91416 379335
rect 90640 379296 90692 379302
rect 90640 379238 90692 379244
rect 91376 379296 91428 379302
rect 91376 379238 91428 379244
rect 92400 379234 92428 379335
rect 92388 379228 92440 379234
rect 92388 379170 92440 379176
rect 90088 378820 90140 378826
rect 90088 378762 90140 378768
rect 86592 378684 86644 378690
rect 86592 378626 86644 378632
rect 93412 378282 93440 380831
rect 110984 380390 111012 380831
rect 110972 380384 111024 380390
rect 110972 380326 111024 380332
rect 113560 380186 113588 380831
rect 116044 380458 116072 380831
rect 118436 380526 118464 380831
rect 118424 380520 118476 380526
rect 118424 380462 118476 380468
rect 116032 380452 116084 380458
rect 116032 380394 116084 380400
rect 121012 380186 121040 380831
rect 123496 380322 123524 380831
rect 123484 380316 123536 380322
rect 123484 380258 123536 380264
rect 125980 380254 126008 380831
rect 131040 380390 131068 380831
rect 133524 380526 133552 380831
rect 133512 380520 133564 380526
rect 133512 380462 133564 380468
rect 135916 380458 135944 380831
rect 146036 380594 146064 380831
rect 146024 380588 146076 380594
rect 146024 380530 146076 380536
rect 135904 380452 135956 380458
rect 135904 380394 135956 380400
rect 131028 380384 131080 380390
rect 128358 380352 128414 380361
rect 131028 380326 131080 380332
rect 155958 380352 156014 380361
rect 128358 380287 128414 380296
rect 155958 380287 156014 380296
rect 128372 380254 128400 380287
rect 125968 380248 126020 380254
rect 125968 380190 126020 380196
rect 128360 380248 128412 380254
rect 128360 380190 128412 380196
rect 113548 380180 113600 380186
rect 113548 380122 113600 380128
rect 121000 380180 121052 380186
rect 121000 380122 121052 380128
rect 155972 380118 156000 380287
rect 155960 380112 156012 380118
rect 155960 380054 156012 380060
rect 158548 380050 158576 380831
rect 160940 380662 160968 380831
rect 160928 380656 160980 380662
rect 160928 380598 160980 380604
rect 163424 380322 163452 380831
rect 163412 380316 163464 380322
rect 163412 380258 163464 380264
rect 158536 380044 158588 380050
rect 158536 379986 158588 379992
rect 166000 379982 166028 380831
rect 165988 379976 166040 379982
rect 165988 379918 166040 379924
rect 93492 379432 93544 379438
rect 93490 379400 93492 379409
rect 93544 379400 93546 379409
rect 93490 379335 93546 379344
rect 96066 379400 96122 379409
rect 96066 379335 96122 379344
rect 98274 379400 98330 379409
rect 98274 379335 98330 379344
rect 98458 379400 98514 379409
rect 98458 379335 98514 379344
rect 101034 379400 101090 379409
rect 101034 379335 101090 379344
rect 103518 379400 103574 379409
rect 103518 379335 103574 379344
rect 105266 379400 105322 379409
rect 105266 379335 105322 379344
rect 108210 379400 108266 379409
rect 108210 379335 108266 379344
rect 108854 379400 108910 379409
rect 108854 379335 108910 379344
rect 111246 379400 111302 379409
rect 111246 379335 111302 379344
rect 112626 379400 112682 379409
rect 112626 379335 112682 379344
rect 113454 379400 113510 379409
rect 113454 379335 113510 379344
rect 114466 379400 114522 379409
rect 114466 379335 114522 379344
rect 117134 379400 117190 379409
rect 117134 379335 117190 379344
rect 141054 379400 141110 379409
rect 141054 379335 141110 379344
rect 148598 379400 148654 379409
rect 148598 379335 148654 379344
rect 150990 379400 151046 379409
rect 150990 379335 151046 379344
rect 153566 379400 153622 379409
rect 153566 379335 153622 379344
rect 183190 379400 183246 379409
rect 183190 379335 183246 379344
rect 95974 379264 96030 379273
rect 95974 379199 96030 379208
rect 94686 378720 94742 378729
rect 94686 378655 94742 378664
rect 93400 378276 93452 378282
rect 93400 378218 93452 378224
rect 85488 378208 85540 378214
rect 85026 378176 85082 378185
rect 85488 378150 85540 378156
rect 85026 378111 85082 378120
rect 83464 376644 83516 376650
rect 83464 376586 83516 376592
rect 85040 375018 85068 378111
rect 94700 376242 94728 378655
rect 94688 376236 94740 376242
rect 94688 376178 94740 376184
rect 95988 376038 96016 379199
rect 96080 378758 96108 379335
rect 96068 378752 96120 378758
rect 96068 378694 96120 378700
rect 97170 378720 97226 378729
rect 97170 378655 97226 378664
rect 97184 376514 97212 378655
rect 98288 377534 98316 379335
rect 98472 379030 98500 379335
rect 99470 379264 99526 379273
rect 99470 379199 99526 379208
rect 98460 379024 98512 379030
rect 98460 378966 98512 378972
rect 98276 377528 98328 377534
rect 98276 377470 98328 377476
rect 97172 376508 97224 376514
rect 97172 376450 97224 376456
rect 99484 376106 99512 379199
rect 101048 378894 101076 379335
rect 102966 379264 103022 379273
rect 102966 379199 103022 379208
rect 101036 378888 101088 378894
rect 101036 378830 101088 378836
rect 101862 378176 101918 378185
rect 101862 378111 101918 378120
rect 99472 376100 99524 376106
rect 99472 376042 99524 376048
rect 95976 376032 96028 376038
rect 95976 375974 96028 375980
rect 101876 375154 101904 378111
rect 102980 375222 103008 379199
rect 103532 378962 103560 379335
rect 105280 379098 105308 379335
rect 105542 379264 105598 379273
rect 105542 379199 105598 379208
rect 105268 379092 105320 379098
rect 105268 379034 105320 379040
rect 103520 378956 103572 378962
rect 103520 378898 103572 378904
rect 104438 378312 104494 378321
rect 104438 378247 104494 378256
rect 104452 375698 104480 378247
rect 105556 377942 105584 379199
rect 108224 379166 108252 379335
rect 108212 379160 108264 379166
rect 108212 379102 108264 379108
rect 108868 378486 108896 379335
rect 108856 378480 108908 378486
rect 108856 378422 108908 378428
rect 111260 378350 111288 379335
rect 112640 379030 112668 379335
rect 112628 379024 112680 379030
rect 112628 378966 112680 378972
rect 113468 378418 113496 379335
rect 114480 379166 114508 379335
rect 114468 379160 114520 379166
rect 114468 379102 114520 379108
rect 117148 379098 117176 379335
rect 117136 379092 117188 379098
rect 117136 379034 117188 379040
rect 138478 378720 138534 378729
rect 138478 378655 138534 378664
rect 113456 378412 113508 378418
rect 113456 378354 113508 378360
rect 111248 378344 111300 378350
rect 107566 378312 107622 378321
rect 111248 378286 111300 378292
rect 107566 378247 107622 378256
rect 106462 378176 106518 378185
rect 106462 378111 106518 378120
rect 105544 377936 105596 377942
rect 105544 377878 105596 377884
rect 104440 375692 104492 375698
rect 104440 375634 104492 375640
rect 106476 375290 106504 378111
rect 107580 375358 107608 378247
rect 138492 376310 138520 378655
rect 141068 377194 141096 379335
rect 148612 377806 148640 379335
rect 151004 377874 151032 379335
rect 150992 377868 151044 377874
rect 150992 377810 151044 377816
rect 148600 377800 148652 377806
rect 148600 377742 148652 377748
rect 153580 377262 153608 379335
rect 182270 378176 182326 378185
rect 182270 378111 182326 378120
rect 182822 378176 182878 378185
rect 182822 378111 182878 378120
rect 182284 378010 182312 378111
rect 182272 378004 182324 378010
rect 182272 377946 182324 377952
rect 153568 377256 153620 377262
rect 153568 377198 153620 377204
rect 141056 377188 141108 377194
rect 141056 377130 141108 377136
rect 138480 376304 138532 376310
rect 138480 376246 138532 376252
rect 107568 375352 107620 375358
rect 107568 375294 107620 375300
rect 106464 375284 106516 375290
rect 106464 375226 106516 375232
rect 102968 375216 103020 375222
rect 102968 375158 103020 375164
rect 101864 375148 101916 375154
rect 101864 375090 101916 375096
rect 85028 375012 85080 375018
rect 85028 374954 85080 374960
rect 178684 360188 178736 360194
rect 178684 360130 178736 360136
rect 178696 358873 178724 360130
rect 179880 360120 179932 360126
rect 179880 360062 179932 360068
rect 179892 358873 179920 360062
rect 178682 358864 178738 358873
rect 178682 358799 178738 358808
rect 179878 358864 179934 358873
rect 179878 358799 179934 358808
rect 182836 358086 182864 378111
rect 183204 378078 183232 379335
rect 183192 378072 183244 378078
rect 183192 378014 183244 378020
rect 196544 360194 196572 381006
rect 196636 377602 196664 488022
rect 196716 484152 196768 484158
rect 196716 484094 196768 484100
rect 196728 377738 196756 484094
rect 196716 377732 196768 377738
rect 196716 377674 196768 377680
rect 196820 377670 196848 488022
rect 196912 488022 197110 488050
rect 196912 484158 196940 488022
rect 197360 485240 197412 485246
rect 197358 485208 197360 485217
rect 197412 485208 197414 485217
rect 197358 485143 197414 485152
rect 197360 485036 197412 485042
rect 197360 484978 197412 484984
rect 197372 484809 197400 484978
rect 197358 484800 197414 484809
rect 197358 484735 197414 484744
rect 197084 484424 197136 484430
rect 197084 484366 197136 484372
rect 196900 484152 196952 484158
rect 196900 484094 196952 484100
rect 196900 471368 196952 471374
rect 196900 471310 196952 471316
rect 196808 377664 196860 377670
rect 196808 377606 196860 377612
rect 196624 377596 196676 377602
rect 196624 377538 196676 377544
rect 196532 360188 196584 360194
rect 196532 360130 196584 360136
rect 196544 359718 196572 360130
rect 196532 359712 196584 359718
rect 196532 359654 196584 359660
rect 190920 359508 190972 359514
rect 190920 359450 190972 359456
rect 190932 358873 190960 359450
rect 190918 358864 190974 358873
rect 190918 358799 190974 358808
rect 60096 358080 60148 358086
rect 60096 358022 60148 358028
rect 182824 358080 182876 358086
rect 182824 358022 182876 358028
rect 95974 273864 96030 273873
rect 95974 273799 96030 273808
rect 113362 273864 113418 273873
rect 113362 273799 113418 273808
rect 76010 273184 76066 273193
rect 76010 273119 76066 273128
rect 77114 273184 77170 273193
rect 77114 273119 77170 273128
rect 90730 273184 90786 273193
rect 90730 273119 90786 273128
rect 93674 273184 93730 273193
rect 93674 273119 93730 273128
rect 94226 273184 94282 273193
rect 94226 273119 94282 273128
rect 60832 272876 60884 272882
rect 60832 272818 60884 272824
rect 60740 272264 60792 272270
rect 60740 272206 60792 272212
rect 60752 252006 60780 272206
rect 60844 272066 60872 272818
rect 76024 272474 76052 273119
rect 77128 272814 77156 273119
rect 77116 272808 77168 272814
rect 77116 272750 77168 272756
rect 90744 272746 90772 273119
rect 90732 272740 90784 272746
rect 90732 272682 90784 272688
rect 93688 272678 93716 273119
rect 94240 272921 94268 273119
rect 94226 272912 94282 272921
rect 94226 272847 94282 272856
rect 94410 272912 94466 272921
rect 94410 272847 94466 272856
rect 95882 272912 95938 272921
rect 95882 272847 95938 272856
rect 93676 272672 93728 272678
rect 93676 272614 93728 272620
rect 76012 272468 76064 272474
rect 76012 272410 76064 272416
rect 94424 272406 94452 272847
rect 95896 272610 95924 272847
rect 95884 272604 95936 272610
rect 95884 272546 95936 272552
rect 62120 272400 62172 272406
rect 94412 272400 94464 272406
rect 62120 272342 62172 272348
rect 83002 272368 83058 272377
rect 60924 272196 60976 272202
rect 60924 272138 60976 272144
rect 60832 272060 60884 272066
rect 60832 272002 60884 272008
rect 60740 252000 60792 252006
rect 60740 251942 60792 251948
rect 60844 251666 60872 272002
rect 60936 252550 60964 272138
rect 62132 271153 62160 272342
rect 94412 272342 94464 272348
rect 83002 272303 83004 272312
rect 83056 272303 83058 272312
rect 83004 272274 83056 272280
rect 95988 272134 96016 273799
rect 98458 272912 98514 272921
rect 98458 272847 98514 272856
rect 98472 272542 98500 272847
rect 98460 272536 98512 272542
rect 98460 272478 98512 272484
rect 107476 272536 107528 272542
rect 107476 272478 107528 272484
rect 100758 272368 100814 272377
rect 100758 272303 100814 272312
rect 100772 272270 100800 272303
rect 100760 272264 100812 272270
rect 99378 272232 99434 272241
rect 100760 272206 100812 272212
rect 99378 272167 99434 272176
rect 102140 272196 102192 272202
rect 95976 272128 96028 272134
rect 95976 272070 96028 272076
rect 98000 271992 98052 271998
rect 98000 271934 98052 271940
rect 98012 271833 98040 271934
rect 84198 271824 84254 271833
rect 84198 271759 84254 271768
rect 97998 271824 98054 271833
rect 97998 271759 98054 271768
rect 62118 271144 62174 271153
rect 62118 271079 62174 271088
rect 61016 270292 61068 270298
rect 61016 270234 61068 270240
rect 81440 270292 81492 270298
rect 81440 270234 81492 270240
rect 61028 269822 61056 270234
rect 80060 269952 80112 269958
rect 80060 269894 80112 269900
rect 61016 269816 61068 269822
rect 61016 269758 61068 269764
rect 60924 252544 60976 252550
rect 60924 252486 60976 252492
rect 61028 252482 61056 269758
rect 80072 268666 80100 269894
rect 80060 268660 80112 268666
rect 80060 268602 80112 268608
rect 81452 268598 81480 270234
rect 84212 269754 84240 271759
rect 88338 271008 88394 271017
rect 88338 270943 88340 270952
rect 88392 270943 88394 270952
rect 89718 271008 89774 271017
rect 89718 270943 89774 270952
rect 88340 270914 88392 270920
rect 85578 270872 85634 270881
rect 85578 270807 85634 270816
rect 88338 270872 88394 270881
rect 88338 270807 88394 270816
rect 84658 270600 84714 270609
rect 84658 270535 84714 270544
rect 84672 270366 84700 270535
rect 84660 270360 84712 270366
rect 84660 270302 84712 270308
rect 85592 270230 85620 270807
rect 86958 270600 87014 270609
rect 86958 270535 87014 270544
rect 86972 270434 87000 270535
rect 86960 270428 87012 270434
rect 86960 270370 87012 270376
rect 88248 270360 88300 270366
rect 88248 270302 88300 270308
rect 85580 270224 85632 270230
rect 85580 270166 85632 270172
rect 86868 270224 86920 270230
rect 86868 270166 86920 270172
rect 84200 269748 84252 269754
rect 84200 269690 84252 269696
rect 81440 268592 81492 268598
rect 81440 268534 81492 268540
rect 86880 268530 86908 270166
rect 86868 268524 86920 268530
rect 86868 268466 86920 268472
rect 88260 268462 88288 270302
rect 88352 270026 88380 270807
rect 89732 270162 89760 270943
rect 92478 270872 92534 270881
rect 92478 270807 92534 270816
rect 91098 270600 91154 270609
rect 91098 270535 91154 270544
rect 89720 270156 89772 270162
rect 89720 270098 89772 270104
rect 88340 270020 88392 270026
rect 88340 269962 88392 269968
rect 91112 269890 91140 270535
rect 92492 270094 92520 270807
rect 92480 270088 92532 270094
rect 92480 270030 92532 270036
rect 91100 269884 91152 269890
rect 91100 269826 91152 269832
rect 88248 268456 88300 268462
rect 88248 268398 88300 268404
rect 99392 268394 99420 272167
rect 102140 272138 102192 272144
rect 102152 271833 102180 272138
rect 104900 272060 104952 272066
rect 104900 272002 104952 272008
rect 104912 271833 104940 272002
rect 107488 271930 107516 272478
rect 107476 271924 107528 271930
rect 107476 271866 107528 271872
rect 107488 271833 107516 271866
rect 102138 271824 102194 271833
rect 102138 271759 102194 271768
rect 104898 271824 104954 271833
rect 104898 271759 104954 271768
rect 107474 271824 107530 271833
rect 107474 271759 107530 271768
rect 100758 271688 100814 271697
rect 100758 271623 100814 271632
rect 110418 271688 110474 271697
rect 110418 271623 110474 271632
rect 100772 271046 100800 271623
rect 103518 271416 103574 271425
rect 103518 271351 103574 271360
rect 103532 271114 103560 271351
rect 110432 271318 110460 271623
rect 113178 271416 113234 271425
rect 113178 271351 113180 271360
rect 113232 271351 113234 271360
rect 113180 271322 113232 271328
rect 110420 271312 110472 271318
rect 104898 271280 104954 271289
rect 104898 271215 104954 271224
rect 107658 271280 107714 271289
rect 110420 271254 110472 271260
rect 107658 271215 107660 271224
rect 104912 271182 104940 271215
rect 107712 271215 107714 271224
rect 107660 271186 107712 271192
rect 104900 271176 104952 271182
rect 104900 271118 104952 271124
rect 111798 271144 111854 271153
rect 103520 271108 103572 271114
rect 111798 271079 111854 271088
rect 103520 271050 103572 271056
rect 100760 271040 100812 271046
rect 100760 270982 100812 270988
rect 106278 270872 106334 270881
rect 106278 270807 106334 270816
rect 99380 268388 99432 268394
rect 99380 268330 99432 268336
rect 61016 252476 61068 252482
rect 61016 252418 61068 252424
rect 106292 251938 106320 270807
rect 109038 270600 109094 270609
rect 109038 270535 109094 270544
rect 110418 270600 110474 270609
rect 110418 270535 110474 270544
rect 109052 270366 109080 270535
rect 109040 270360 109092 270366
rect 109040 270302 109092 270308
rect 110432 270230 110460 270535
rect 111812 270298 111840 271079
rect 111800 270292 111852 270298
rect 111800 270234 111852 270240
rect 110420 270224 110472 270230
rect 110420 270166 110472 270172
rect 113376 269890 113404 273799
rect 133418 273728 133474 273737
rect 133418 273663 133474 273672
rect 133432 273630 133460 273663
rect 133420 273624 133472 273630
rect 133420 273566 133472 273572
rect 135902 273592 135958 273601
rect 135902 273527 135904 273536
rect 135956 273527 135958 273536
rect 138478 273592 138534 273601
rect 138478 273527 138534 273536
rect 140870 273592 140926 273601
rect 140870 273527 140926 273536
rect 143538 273592 143594 273601
rect 143538 273527 143594 273536
rect 145930 273592 145986 273601
rect 145930 273527 145986 273536
rect 135904 273498 135956 273504
rect 138492 273494 138520 273527
rect 138480 273488 138532 273494
rect 138480 273430 138532 273436
rect 140884 273426 140912 273527
rect 140872 273420 140924 273426
rect 140872 273362 140924 273368
rect 143552 273358 143580 273527
rect 143540 273352 143592 273358
rect 143540 273294 143592 273300
rect 145944 273290 145972 273527
rect 145932 273284 145984 273290
rect 145932 273226 145984 273232
rect 196912 272542 196940 471310
rect 196992 380996 197044 381002
rect 196992 380938 197044 380944
rect 196900 272536 196952 272542
rect 196900 272478 196952 272484
rect 114468 271924 114520 271930
rect 114468 271866 114520 271872
rect 127624 271924 127676 271930
rect 127624 271866 127676 271872
rect 114480 271833 114508 271866
rect 114466 271824 114522 271833
rect 114466 271759 114522 271768
rect 123206 271824 123262 271833
rect 123206 271759 123208 271768
rect 123260 271759 123262 271768
rect 125598 271824 125654 271833
rect 125598 271759 125654 271768
rect 123208 271730 123260 271736
rect 125612 271726 125640 271759
rect 125600 271720 125652 271726
rect 120078 271688 120134 271697
rect 125600 271662 125652 271668
rect 120078 271623 120134 271632
rect 120092 271590 120120 271623
rect 120080 271584 120132 271590
rect 115938 271552 115994 271561
rect 115938 271487 115940 271496
rect 115992 271487 115994 271496
rect 117318 271552 117374 271561
rect 120080 271526 120132 271532
rect 117318 271487 117374 271496
rect 115940 271458 115992 271464
rect 117332 271454 117360 271487
rect 117320 271448 117372 271454
rect 117320 271390 117372 271396
rect 118698 271280 118754 271289
rect 118698 271215 118754 271224
rect 114558 271008 114614 271017
rect 114558 270943 114614 270952
rect 114572 269958 114600 270943
rect 115938 270872 115994 270881
rect 115938 270807 115994 270816
rect 114560 269952 114612 269958
rect 114560 269894 114612 269900
rect 113364 269884 113416 269890
rect 113364 269826 113416 269832
rect 106280 251932 106332 251938
rect 106280 251874 106332 251880
rect 115952 251870 115980 270807
rect 118712 269822 118740 271215
rect 127636 271182 127664 271866
rect 129740 271856 129792 271862
rect 129738 271824 129740 271833
rect 154488 271856 154540 271862
rect 129792 271824 129794 271833
rect 129738 271759 129794 271768
rect 151358 271824 151414 271833
rect 151358 271759 151414 271768
rect 154486 271824 154488 271833
rect 154540 271824 154542 271833
rect 154486 271759 154542 271768
rect 158626 271824 158682 271833
rect 158626 271759 158628 271768
rect 151372 271726 151400 271759
rect 158680 271759 158682 271768
rect 158628 271730 158680 271736
rect 151360 271720 151412 271726
rect 128358 271688 128414 271697
rect 151360 271662 151412 271668
rect 157246 271688 157302 271697
rect 128358 271623 128360 271632
rect 128412 271623 128414 271632
rect 157246 271623 157248 271632
rect 128360 271594 128412 271600
rect 157300 271623 157302 271632
rect 161294 271688 161350 271697
rect 161294 271623 161350 271632
rect 164146 271688 164202 271697
rect 164146 271623 164202 271632
rect 166906 271688 166962 271697
rect 166906 271623 166962 271632
rect 183466 271688 183522 271697
rect 183466 271623 183522 271632
rect 157248 271594 157300 271600
rect 161308 271590 161336 271623
rect 161296 271584 161348 271590
rect 161296 271526 161348 271532
rect 164160 271522 164188 271623
rect 164148 271516 164200 271522
rect 164148 271458 164200 271464
rect 166920 271454 166948 271623
rect 166908 271448 166960 271454
rect 166908 271390 166960 271396
rect 183480 271250 183508 271623
rect 196624 271448 196676 271454
rect 196624 271390 196676 271396
rect 183468 271244 183520 271250
rect 183468 271186 183520 271192
rect 196636 271182 196664 271390
rect 127624 271176 127676 271182
rect 127624 271118 127676 271124
rect 196624 271176 196676 271182
rect 196624 271118 196676 271124
rect 147678 270872 147734 270881
rect 147678 270807 147734 270816
rect 147692 270502 147720 270807
rect 183466 270600 183522 270609
rect 183466 270535 183468 270544
rect 183520 270535 183522 270544
rect 183468 270506 183520 270512
rect 147680 270496 147732 270502
rect 147680 270438 147732 270444
rect 128360 269884 128412 269890
rect 128360 269826 128412 269832
rect 118700 269816 118752 269822
rect 118700 269758 118752 269764
rect 128372 269074 128400 269826
rect 128360 269068 128412 269074
rect 128360 269010 128412 269016
rect 180156 253360 180208 253366
rect 180154 253328 180156 253337
rect 180208 253328 180210 253337
rect 179328 253292 179380 253298
rect 180154 253263 180210 253272
rect 179328 253234 179380 253240
rect 179340 253201 179368 253234
rect 191748 253224 191800 253230
rect 179326 253192 179382 253201
rect 179326 253127 179382 253136
rect 191746 253192 191748 253201
rect 191800 253192 191802 253201
rect 191746 253127 191802 253136
rect 115940 251864 115992 251870
rect 115940 251806 115992 251812
rect 60832 251660 60884 251666
rect 60832 251602 60884 251608
rect 96068 167000 96120 167006
rect 96068 166942 96120 166948
rect 96080 166841 96108 166942
rect 98460 166932 98512 166938
rect 98460 166874 98512 166880
rect 98472 166841 98500 166874
rect 101036 166864 101088 166870
rect 96066 166832 96122 166841
rect 96066 166767 96122 166776
rect 98458 166832 98514 166841
rect 98458 166767 98514 166776
rect 101034 166832 101036 166841
rect 101088 166832 101090 166841
rect 101034 166767 101090 166776
rect 105818 166832 105874 166841
rect 105818 166767 105820 166776
rect 105872 166767 105874 166776
rect 108210 166832 108266 166841
rect 108210 166767 108266 166776
rect 138478 166832 138534 166841
rect 138478 166767 138534 166776
rect 140870 166832 140926 166841
rect 140870 166767 140926 166776
rect 145930 166832 145986 166841
rect 145930 166767 145986 166776
rect 105820 166738 105872 166744
rect 108224 166734 108252 166767
rect 108212 166728 108264 166734
rect 108212 166670 108264 166676
rect 138492 166598 138520 166767
rect 140884 166666 140912 166767
rect 140872 166660 140924 166666
rect 140872 166602 140924 166608
rect 138480 166592 138532 166598
rect 111154 166560 111210 166569
rect 111154 166495 111210 166504
rect 116950 166560 117006 166569
rect 138480 166534 138532 166540
rect 145944 166530 145972 166767
rect 163318 166696 163374 166705
rect 163318 166631 163374 166640
rect 148506 166560 148562 166569
rect 116950 166495 117006 166504
rect 145932 166524 145984 166530
rect 60740 166252 60792 166258
rect 60740 166194 60792 166200
rect 60752 146130 60780 166194
rect 111168 165714 111196 166495
rect 111156 165708 111208 165714
rect 111156 165650 111208 165656
rect 116964 165646 116992 166495
rect 148506 166495 148562 166504
rect 145932 166466 145984 166472
rect 148520 166462 148548 166495
rect 148508 166456 148560 166462
rect 148508 166398 148560 166404
rect 153290 166424 153346 166433
rect 153290 166359 153292 166368
rect 153344 166359 153346 166368
rect 153292 166330 153344 166336
rect 163332 166326 163360 166631
rect 163320 166320 163372 166326
rect 163320 166262 163372 166268
rect 116952 165640 117004 165646
rect 81438 165608 81494 165617
rect 81438 165543 81494 165552
rect 84198 165608 84254 165617
rect 84198 165543 84254 165552
rect 91190 165608 91246 165617
rect 91190 165543 91246 165552
rect 95238 165608 95294 165617
rect 95238 165543 95294 165552
rect 99378 165608 99434 165617
rect 99378 165543 99434 165552
rect 103518 165608 103574 165617
rect 103518 165543 103574 165552
rect 109314 165608 109370 165617
rect 109314 165543 109370 165552
rect 110970 165608 111026 165617
rect 110970 165543 111026 165552
rect 113546 165608 113602 165617
rect 113546 165543 113602 165552
rect 115938 165608 115994 165617
rect 116952 165582 117004 165588
rect 117870 165608 117926 165617
rect 115938 165543 115994 165552
rect 117870 165543 117926 165552
rect 118146 165608 118202 165617
rect 118146 165543 118202 165552
rect 120906 165608 120962 165617
rect 120906 165543 120962 165552
rect 123482 165608 123538 165617
rect 123482 165543 123538 165552
rect 125874 165608 125930 165617
rect 125874 165543 125930 165552
rect 128358 165608 128414 165617
rect 128358 165543 128414 165552
rect 129738 165608 129794 165617
rect 129738 165543 129794 165552
rect 132498 165608 132554 165617
rect 132498 165543 132554 165552
rect 135258 165608 135314 165617
rect 135258 165543 135314 165552
rect 150438 165608 150494 165617
rect 150438 165543 150440 165552
rect 75918 164384 75974 164393
rect 75918 164319 75974 164328
rect 60740 146124 60792 146130
rect 60740 146066 60792 146072
rect 66260 146124 66312 146130
rect 66260 146066 66312 146072
rect 66272 146010 66300 146066
rect 66444 146056 66496 146062
rect 66272 146004 66444 146010
rect 66272 145998 66496 146004
rect 66272 145982 66484 145998
rect 75932 145450 75960 164319
rect 76010 164248 76066 164257
rect 76010 164183 76066 164192
rect 77298 164248 77354 164257
rect 77298 164183 77354 164192
rect 78678 164248 78734 164257
rect 78678 164183 78734 164192
rect 80058 164248 80114 164257
rect 80058 164183 80114 164192
rect 75920 145444 75972 145450
rect 75920 145386 75972 145392
rect 76024 145382 76052 164183
rect 77312 145518 77340 164183
rect 78692 148782 78720 164183
rect 80072 148850 80100 164183
rect 80060 148844 80112 148850
rect 80060 148786 80112 148792
rect 78680 148776 78732 148782
rect 78680 148718 78732 148724
rect 81452 148714 81480 165543
rect 82818 164248 82874 164257
rect 82818 164183 82874 164192
rect 81440 148708 81492 148714
rect 81440 148650 81492 148656
rect 82832 145654 82860 164183
rect 84212 145790 84240 165543
rect 88338 164792 88394 164801
rect 88338 164727 88394 164736
rect 89994 164792 90050 164801
rect 89994 164727 89996 164736
rect 88352 164694 88380 164727
rect 90048 164727 90050 164736
rect 89996 164698 90048 164704
rect 88340 164688 88392 164694
rect 88340 164630 88392 164636
rect 84290 164248 84346 164257
rect 84290 164183 84346 164192
rect 85578 164248 85634 164257
rect 85578 164183 85634 164192
rect 86958 164248 87014 164257
rect 86958 164183 87014 164192
rect 88430 164248 88486 164257
rect 88430 164183 88486 164192
rect 89810 164248 89866 164257
rect 89810 164183 89866 164192
rect 91098 164248 91154 164257
rect 91098 164183 91154 164192
rect 84200 145784 84252 145790
rect 84200 145726 84252 145732
rect 84304 145722 84332 164183
rect 85592 145858 85620 164183
rect 86972 146198 87000 164183
rect 86960 146192 87012 146198
rect 86960 146134 87012 146140
rect 88444 145994 88472 164183
rect 88432 145988 88484 145994
rect 88432 145930 88484 145936
rect 89824 145926 89852 164183
rect 91112 146266 91140 164183
rect 91100 146260 91152 146266
rect 91100 146202 91152 146208
rect 89812 145920 89864 145926
rect 89812 145862 89864 145868
rect 85580 145852 85632 145858
rect 85580 145794 85632 145800
rect 84292 145716 84344 145722
rect 84292 145658 84344 145664
rect 82820 145648 82872 145654
rect 82820 145590 82872 145596
rect 91204 145586 91232 165543
rect 91744 164892 91796 164898
rect 91744 164834 91796 164840
rect 91756 164694 91784 164834
rect 94596 164824 94648 164830
rect 94780 164824 94832 164830
rect 94648 164772 94780 164778
rect 94596 164766 94832 164772
rect 94608 164750 94820 164766
rect 91744 164688 91796 164694
rect 91744 164630 91796 164636
rect 92478 164248 92534 164257
rect 92478 164183 92534 164192
rect 93858 164248 93914 164257
rect 93858 164183 93914 164192
rect 92492 146130 92520 164183
rect 92480 146124 92532 146130
rect 92480 146066 92532 146072
rect 93872 146062 93900 164183
rect 95252 163878 95280 165543
rect 96618 164520 96674 164529
rect 96618 164455 96674 164464
rect 95240 163872 95292 163878
rect 95240 163814 95292 163820
rect 96632 163810 96660 164455
rect 98644 164348 98696 164354
rect 98644 164290 98696 164296
rect 97998 164248 98054 164257
rect 97998 164183 98054 164192
rect 96620 163804 96672 163810
rect 96620 163746 96672 163752
rect 98012 163742 98040 164183
rect 98000 163736 98052 163742
rect 98000 163678 98052 163684
rect 93860 146056 93912 146062
rect 93860 145998 93912 146004
rect 98656 145625 98684 164290
rect 99392 145761 99420 165543
rect 103532 164694 103560 165543
rect 103520 164688 103572 164694
rect 103520 164630 103572 164636
rect 100758 164384 100814 164393
rect 100758 164319 100760 164328
rect 100812 164319 100814 164328
rect 103518 164384 103574 164393
rect 103518 164319 103574 164328
rect 100760 164290 100812 164296
rect 103532 164286 103560 164319
rect 100024 164280 100076 164286
rect 103520 164280 103572 164286
rect 100024 164222 100076 164228
rect 100758 164248 100814 164257
rect 100036 148646 100064 164222
rect 100758 164183 100814 164192
rect 102138 164248 102194 164257
rect 103520 164222 103572 164228
rect 106186 164248 106242 164257
rect 102138 164183 102194 164192
rect 106370 164248 106426 164257
rect 106242 164206 106320 164234
rect 106186 164183 106242 164192
rect 100024 148640 100076 148646
rect 100024 148582 100076 148588
rect 100772 145897 100800 164183
rect 102152 146305 102180 164183
rect 106292 149054 106320 164206
rect 106370 164183 106426 164192
rect 107566 164248 107622 164257
rect 107622 164206 107792 164234
rect 107566 164183 107622 164192
rect 106384 163674 106412 164183
rect 107658 164112 107714 164121
rect 107658 164047 107714 164056
rect 106372 163668 106424 163674
rect 106372 163610 106424 163616
rect 106280 149048 106332 149054
rect 106280 148990 106332 148996
rect 107672 148578 107700 164047
rect 107660 148572 107712 148578
rect 107660 148514 107712 148520
rect 107764 148510 107792 164206
rect 109328 163606 109356 165543
rect 110984 164150 111012 165543
rect 113560 164966 113588 165543
rect 115952 165034 115980 165543
rect 115940 165028 115992 165034
rect 115940 164970 115992 164976
rect 113548 164960 113600 164966
rect 114652 164960 114704 164966
rect 113548 164902 113600 164908
rect 114466 164928 114522 164937
rect 114652 164902 114704 164908
rect 114466 164863 114468 164872
rect 114520 164863 114522 164872
rect 114468 164834 114520 164840
rect 112074 164656 112130 164665
rect 112074 164591 112130 164600
rect 110972 164144 111024 164150
rect 110972 164086 111024 164092
rect 109316 163600 109368 163606
rect 109316 163542 109368 163548
rect 112088 162246 112116 164591
rect 114664 164529 114692 164902
rect 114744 164892 114796 164898
rect 114744 164834 114796 164840
rect 114650 164520 114706 164529
rect 114650 164455 114706 164464
rect 112076 162240 112128 162246
rect 112076 162182 112128 162188
rect 107752 148504 107804 148510
rect 107752 148446 107804 148452
rect 114664 148442 114692 164455
rect 114652 148436 114704 148442
rect 114652 148378 114704 148384
rect 114756 148374 114784 164834
rect 115754 164656 115810 164665
rect 115754 164591 115810 164600
rect 115768 162178 115796 164591
rect 117884 164218 117912 165543
rect 118160 164830 118188 165543
rect 120920 165102 120948 165543
rect 123496 165170 123524 165543
rect 125888 165238 125916 165543
rect 128372 165374 128400 165543
rect 128360 165368 128412 165374
rect 128360 165310 128412 165316
rect 129752 165306 129780 165543
rect 132512 165442 132540 165543
rect 135272 165510 135300 165543
rect 150492 165543 150494 165552
rect 183190 165608 183246 165617
rect 183190 165543 183246 165552
rect 183466 165608 183522 165617
rect 183466 165543 183522 165552
rect 150440 165514 150492 165520
rect 135260 165504 135312 165510
rect 135260 165446 135312 165452
rect 132500 165436 132552 165442
rect 132500 165378 132552 165384
rect 129740 165300 129792 165306
rect 129740 165242 129792 165248
rect 125876 165232 125928 165238
rect 125876 165174 125928 165180
rect 123484 165164 123536 165170
rect 123484 165106 123536 165112
rect 120908 165096 120960 165102
rect 118882 165064 118938 165073
rect 120908 165038 120960 165044
rect 183204 165034 183232 165543
rect 183480 165170 183508 165543
rect 183468 165164 183520 165170
rect 183468 165106 183520 165112
rect 118882 164999 118938 165008
rect 183192 165028 183244 165034
rect 118148 164824 118200 164830
rect 118148 164766 118200 164772
rect 117872 164212 117924 164218
rect 117872 164154 117924 164160
rect 118896 163538 118924 164999
rect 183192 164970 183244 164976
rect 196636 164898 196664 271118
rect 197004 269074 197032 380938
rect 197096 377398 197124 484366
rect 197452 484152 197504 484158
rect 197452 484094 197504 484100
rect 197176 482588 197228 482594
rect 197176 482530 197228 482536
rect 197188 465050 197216 482530
rect 197268 468716 197320 468722
rect 197268 468658 197320 468664
rect 197176 465044 197228 465050
rect 197176 464986 197228 464992
rect 197176 381540 197228 381546
rect 197176 381482 197228 381488
rect 197084 377392 197136 377398
rect 197084 377334 197136 377340
rect 197188 373994 197216 381482
rect 197280 377806 197308 468658
rect 197464 378010 197492 484094
rect 197452 378004 197504 378010
rect 197452 377946 197504 377952
rect 197556 377806 197584 488036
rect 198046 488022 198320 488050
rect 197912 482520 197964 482526
rect 197912 482462 197964 482468
rect 197728 468648 197780 468654
rect 197728 468590 197780 468596
rect 197636 468580 197688 468586
rect 197636 468522 197688 468528
rect 197268 377800 197320 377806
rect 197268 377742 197320 377748
rect 197544 377800 197596 377806
rect 197544 377742 197596 377748
rect 197188 373966 197308 373994
rect 197280 360126 197308 373966
rect 197268 360120 197320 360126
rect 197268 360062 197320 360068
rect 197280 359802 197308 360062
rect 197280 359774 197492 359802
rect 197360 359712 197412 359718
rect 197360 359654 197412 359660
rect 196992 269068 197044 269074
rect 196992 269010 197044 269016
rect 197004 258074 197032 269010
rect 196728 258046 197032 258074
rect 196728 164966 196756 258046
rect 197372 253298 197400 359654
rect 197464 354674 197492 359774
rect 197464 354646 197584 354674
rect 197452 271244 197504 271250
rect 197452 271186 197504 271192
rect 197360 253292 197412 253298
rect 197360 253234 197412 253240
rect 197360 165572 197412 165578
rect 197360 165514 197412 165520
rect 197372 165170 197400 165514
rect 197360 165164 197412 165170
rect 197360 165106 197412 165112
rect 196716 164960 196768 164966
rect 196716 164902 196768 164908
rect 196624 164892 196676 164898
rect 196624 164834 196676 164840
rect 118884 163532 118936 163538
rect 118884 163474 118936 163480
rect 115756 162172 115808 162178
rect 115756 162114 115808 162120
rect 114744 148368 114796 148374
rect 114744 148310 114796 148316
rect 102138 146296 102194 146305
rect 102138 146231 102194 146240
rect 179052 146260 179104 146266
rect 179052 146202 179104 146208
rect 100758 145888 100814 145897
rect 100758 145823 100814 145832
rect 99378 145752 99434 145761
rect 99378 145687 99434 145696
rect 98642 145616 98698 145625
rect 91192 145580 91244 145586
rect 98642 145551 98698 145560
rect 91192 145522 91244 145528
rect 77300 145512 77352 145518
rect 77300 145454 77352 145460
rect 76012 145376 76064 145382
rect 76012 145318 76064 145324
rect 179064 144945 179092 146202
rect 179696 146192 179748 146198
rect 179696 146134 179748 146140
rect 179708 144945 179736 146134
rect 191288 145580 191340 145586
rect 191288 145522 191340 145528
rect 191300 144945 191328 145522
rect 179050 144936 179106 144945
rect 179050 144871 179106 144880
rect 179694 144936 179750 144945
rect 179694 144871 179750 144880
rect 191286 144936 191342 144945
rect 191286 144871 191342 144880
rect 77114 59800 77170 59809
rect 77114 59735 77116 59744
rect 77168 59735 77170 59744
rect 83094 59800 83150 59809
rect 83094 59735 83150 59744
rect 101770 59800 101826 59809
rect 101770 59735 101826 59744
rect 103886 59800 103942 59809
rect 103886 59735 103942 59744
rect 107566 59800 107622 59809
rect 107566 59735 107622 59744
rect 113546 59800 113602 59809
rect 113546 59735 113602 59744
rect 77116 59706 77168 59712
rect 83108 59702 83136 59735
rect 83096 59696 83148 59702
rect 83096 59638 83148 59644
rect 94502 59664 94558 59673
rect 94502 59599 94558 59608
rect 96986 59664 97042 59673
rect 96986 59599 97042 59608
rect 98090 59664 98146 59673
rect 98090 59599 98146 59608
rect 100758 59664 100814 59673
rect 100758 59599 100760 59608
rect 84200 59356 84252 59362
rect 84200 59298 84252 59304
rect 84212 58041 84240 59298
rect 94516 59294 94544 59599
rect 95882 59528 95938 59537
rect 95882 59463 95938 59472
rect 94504 59288 94556 59294
rect 94504 59230 94556 59236
rect 95896 59226 95924 59463
rect 95884 59220 95936 59226
rect 95884 59162 95936 59168
rect 97000 59158 97028 59599
rect 96988 59152 97040 59158
rect 96988 59094 97040 59100
rect 98104 59090 98132 59599
rect 100812 59599 100814 59608
rect 100760 59570 100812 59576
rect 101784 59566 101812 59735
rect 102782 59664 102838 59673
rect 102782 59599 102838 59608
rect 101772 59560 101824 59566
rect 101772 59502 101824 59508
rect 98092 59084 98144 59090
rect 98092 59026 98144 59032
rect 102796 59022 102824 59599
rect 102784 59016 102836 59022
rect 102784 58958 102836 58964
rect 103900 58954 103928 59735
rect 107580 59498 107608 59735
rect 108670 59664 108726 59673
rect 108670 59599 108726 59608
rect 107568 59492 107620 59498
rect 107568 59434 107620 59440
rect 103888 58948 103940 58954
rect 103888 58890 103940 58896
rect 108684 58886 108712 59599
rect 113560 59430 113588 59735
rect 113548 59424 113600 59430
rect 110970 59392 111026 59401
rect 113548 59366 113600 59372
rect 110970 59327 111026 59336
rect 108672 58880 108724 58886
rect 108672 58822 108724 58828
rect 110984 58818 111012 59327
rect 148506 59256 148562 59265
rect 148506 59191 148562 59200
rect 150898 59256 150954 59265
rect 150898 59191 150954 59200
rect 110972 58812 111024 58818
rect 110972 58754 111024 58760
rect 148520 58750 148548 59191
rect 148508 58744 148560 58750
rect 148508 58686 148560 58692
rect 150912 58682 150940 59191
rect 150900 58676 150952 58682
rect 150900 58618 150952 58624
rect 84198 58032 84254 58041
rect 84198 57967 84254 57976
rect 76010 57896 76066 57905
rect 76010 57831 76066 57840
rect 78218 57896 78274 57905
rect 78218 57831 78274 57840
rect 79506 57896 79562 57905
rect 79506 57831 79562 57840
rect 80058 57896 80114 57905
rect 80058 57831 80114 57840
rect 81898 57896 81954 57905
rect 81898 57831 81954 57840
rect 85394 57896 85450 57905
rect 85394 57831 85450 57840
rect 86498 57896 86554 57905
rect 86498 57831 86554 57840
rect 86958 57896 87014 57905
rect 86958 57831 87014 57840
rect 88706 57896 88762 57905
rect 88706 57831 88762 57840
rect 89810 57896 89866 57905
rect 89810 57831 89866 57840
rect 90730 57896 90786 57905
rect 90730 57831 90786 57840
rect 91190 57896 91246 57905
rect 91190 57831 91246 57840
rect 92202 57896 92258 57905
rect 92202 57831 92258 57840
rect 92478 57896 92534 57905
rect 92478 57831 92534 57840
rect 93582 57896 93638 57905
rect 93582 57831 93638 57840
rect 99378 57896 99434 57905
rect 99378 57831 99434 57840
rect 109498 57896 109554 57905
rect 109498 57831 109554 57840
rect 112074 57896 112130 57905
rect 112074 57831 112130 57840
rect 113822 57896 113878 57905
rect 113822 57831 113878 57840
rect 115938 57896 115994 57905
rect 115938 57831 115994 57840
rect 116674 57896 116730 57905
rect 116674 57831 116730 57840
rect 123482 57896 123538 57905
rect 123482 57831 123538 57840
rect 125874 57896 125930 57905
rect 125874 57831 125930 57840
rect 128358 57896 128414 57905
rect 128358 57831 128414 57840
rect 130842 57896 130898 57905
rect 130842 57831 130898 57840
rect 133418 57896 133474 57905
rect 133418 57831 133474 57840
rect 145562 57896 145618 57905
rect 145562 57831 145564 57840
rect 60004 57452 60056 57458
rect 60004 57394 60056 57400
rect 76024 57186 76052 57831
rect 78232 57254 78260 57831
rect 78220 57248 78272 57254
rect 78220 57190 78272 57196
rect 76012 57180 76064 57186
rect 76012 57122 76064 57128
rect 79520 55894 79548 57831
rect 79508 55888 79560 55894
rect 79508 55830 79560 55836
rect 59912 55004 59964 55010
rect 59912 54946 59964 54952
rect 59176 54732 59228 54738
rect 59176 54674 59228 54680
rect 80072 54670 80100 57831
rect 81912 56030 81940 57831
rect 81900 56024 81952 56030
rect 81900 55966 81952 55972
rect 85408 55962 85436 57831
rect 86512 56098 86540 57831
rect 86500 56092 86552 56098
rect 86500 56034 86552 56040
rect 85396 55956 85448 55962
rect 85396 55898 85448 55904
rect 86972 54874 87000 57831
rect 88720 56166 88748 57831
rect 88708 56160 88760 56166
rect 88708 56102 88760 56108
rect 86960 54868 87012 54874
rect 86960 54810 87012 54816
rect 89824 54738 89852 57831
rect 90744 56302 90772 57831
rect 90732 56296 90784 56302
rect 90732 56238 90784 56244
rect 91204 54942 91232 57831
rect 92216 56234 92244 57831
rect 92204 56228 92256 56234
rect 92204 56170 92256 56176
rect 91192 54936 91244 54942
rect 91192 54878 91244 54884
rect 92492 54806 92520 57831
rect 93596 57322 93624 57831
rect 98550 57488 98606 57497
rect 98550 57423 98606 57432
rect 93584 57316 93636 57322
rect 93584 57258 93636 57264
rect 98564 57225 98592 57423
rect 99392 57390 99420 57831
rect 106278 57624 106334 57633
rect 106278 57559 106334 57568
rect 99380 57384 99432 57390
rect 99380 57326 99432 57332
rect 98550 57216 98606 57225
rect 98550 57151 98606 57160
rect 106292 55010 106320 57559
rect 109512 56370 109540 57831
rect 110418 57624 110474 57633
rect 110418 57559 110474 57568
rect 109500 56364 109552 56370
rect 109500 56306 109552 56312
rect 110432 55078 110460 57559
rect 112088 56438 112116 57831
rect 113270 57624 113326 57633
rect 113270 57559 113326 57568
rect 112076 56432 112128 56438
rect 112076 56374 112128 56380
rect 113284 55146 113312 57559
rect 113836 56506 113864 57831
rect 114558 57624 114614 57633
rect 114558 57559 114614 57568
rect 113824 56500 113876 56506
rect 113824 56442 113876 56448
rect 114572 55214 114600 57559
rect 115952 57526 115980 57831
rect 115940 57520 115992 57526
rect 115940 57462 115992 57468
rect 116688 56574 116716 57831
rect 123496 57798 123524 57831
rect 123484 57792 123536 57798
rect 123484 57734 123536 57740
rect 118698 57624 118754 57633
rect 118698 57559 118754 57568
rect 116676 56568 116728 56574
rect 116676 56510 116728 56516
rect 114560 55208 114612 55214
rect 114560 55150 114612 55156
rect 113272 55140 113324 55146
rect 113272 55082 113324 55088
rect 110420 55072 110472 55078
rect 110420 55014 110472 55020
rect 106280 55004 106332 55010
rect 106280 54946 106332 54952
rect 92480 54800 92532 54806
rect 118712 54777 118740 57559
rect 125888 57458 125916 57831
rect 128372 57594 128400 57831
rect 130856 57662 130884 57831
rect 133432 57730 133460 57831
rect 145616 57831 145618 57840
rect 153290 57896 153346 57905
rect 153290 57831 153346 57840
rect 183282 57896 183338 57905
rect 183282 57831 183284 57840
rect 145564 57802 145616 57808
rect 133420 57724 133472 57730
rect 133420 57666 133472 57672
rect 130844 57656 130896 57662
rect 130844 57598 130896 57604
rect 128360 57588 128412 57594
rect 128360 57530 128412 57536
rect 125876 57452 125928 57458
rect 125876 57394 125928 57400
rect 153304 56273 153332 57831
rect 183336 57831 183338 57840
rect 183284 57802 183336 57808
rect 197372 57798 197400 165106
rect 197464 165034 197492 271186
rect 197556 253366 197584 354646
rect 197648 271726 197676 468522
rect 197636 271720 197688 271726
rect 197636 271662 197688 271668
rect 197740 271522 197768 468590
rect 197820 464500 197872 464506
rect 197820 464442 197872 464448
rect 197728 271516 197780 271522
rect 197728 271458 197780 271464
rect 197832 271454 197860 464442
rect 197924 380186 197952 482462
rect 198004 464432 198056 464438
rect 198004 464374 198056 464380
rect 198016 380322 198044 464374
rect 198186 398032 198242 398041
rect 198186 397967 198242 397976
rect 198096 397860 198148 397866
rect 198096 397802 198148 397808
rect 198004 380316 198056 380322
rect 198004 380258 198056 380264
rect 197912 380180 197964 380186
rect 197912 380122 197964 380128
rect 198004 378072 198056 378078
rect 198004 378014 198056 378020
rect 198016 374950 198044 378014
rect 198108 377874 198136 397802
rect 198200 381002 198228 397967
rect 198188 380996 198240 381002
rect 198188 380938 198240 380944
rect 198292 377874 198320 488022
rect 198384 488022 198490 488050
rect 198384 484158 198412 488022
rect 198372 484152 198424 484158
rect 198372 484094 198424 484100
rect 198740 484152 198792 484158
rect 198740 484094 198792 484100
rect 198096 377868 198148 377874
rect 198096 377810 198148 377816
rect 198280 377868 198332 377874
rect 198280 377810 198332 377816
rect 198752 377330 198780 484094
rect 198844 378078 198872 488036
rect 198936 488022 199318 488050
rect 199794 488022 199884 488050
rect 198936 484158 198964 488022
rect 199108 486532 199160 486538
rect 199108 486474 199160 486480
rect 198924 484152 198976 484158
rect 198924 484094 198976 484100
rect 199016 468784 199068 468790
rect 199016 468726 199068 468732
rect 198924 465724 198976 465730
rect 198924 465666 198976 465672
rect 198936 465118 198964 465666
rect 198924 465112 198976 465118
rect 198924 465054 198976 465060
rect 198936 460193 198964 465054
rect 198922 460184 198978 460193
rect 198922 460119 198978 460128
rect 198832 378072 198884 378078
rect 198832 378014 198884 378020
rect 198740 377324 198792 377330
rect 198740 377266 198792 377272
rect 198004 374944 198056 374950
rect 198004 374886 198056 374892
rect 197820 271448 197872 271454
rect 197820 271390 197872 271396
rect 197912 271312 197964 271318
rect 197912 271254 197964 271260
rect 197924 270570 197952 271254
rect 198016 271250 198044 374886
rect 198936 354674 198964 460119
rect 199028 379982 199056 468726
rect 199120 397866 199148 486474
rect 199384 485308 199436 485314
rect 199384 485250 199436 485256
rect 199200 479528 199252 479534
rect 199200 479470 199252 479476
rect 199212 398274 199240 479470
rect 199292 464364 199344 464370
rect 199292 464306 199344 464312
rect 199200 398268 199252 398274
rect 199200 398210 199252 398216
rect 199198 398168 199254 398177
rect 199198 398103 199254 398112
rect 199108 397860 199160 397866
rect 199108 397802 199160 397808
rect 199106 396808 199162 396817
rect 199106 396743 199162 396752
rect 199016 379976 199068 379982
rect 199016 379918 199068 379924
rect 199014 379400 199070 379409
rect 199014 379335 199070 379344
rect 199028 378826 199056 379335
rect 199016 378820 199068 378826
rect 199016 378762 199068 378768
rect 199028 378622 199056 378762
rect 199016 378616 199068 378622
rect 199016 378558 199068 378564
rect 199120 378146 199148 396743
rect 199212 396137 199240 398103
rect 199198 396128 199254 396137
rect 199198 396063 199254 396072
rect 199304 380254 199332 464306
rect 199292 380248 199344 380254
rect 199292 380190 199344 380196
rect 199108 378140 199160 378146
rect 199108 378082 199160 378088
rect 199396 377466 199424 485250
rect 199856 485246 199884 488022
rect 200224 485353 200252 488036
rect 200316 488022 200698 488050
rect 200776 488022 201066 488050
rect 201542 488022 201632 488050
rect 200210 485344 200266 485353
rect 200210 485279 200266 485288
rect 199844 485240 199896 485246
rect 199844 485182 199896 485188
rect 200316 484106 200344 488022
rect 200488 484900 200540 484906
rect 200488 484842 200540 484848
rect 200500 484809 200528 484842
rect 200486 484800 200542 484809
rect 200486 484735 200542 484744
rect 200132 484078 200344 484106
rect 199568 475380 199620 475386
rect 199568 475322 199620 475328
rect 199476 465656 199528 465662
rect 199476 465598 199528 465604
rect 199488 381002 199516 465598
rect 199580 400353 199608 475322
rect 199566 400344 199622 400353
rect 199566 400279 199622 400288
rect 199476 380996 199528 381002
rect 199476 380938 199528 380944
rect 199474 377904 199530 377913
rect 199474 377839 199530 377848
rect 199384 377460 199436 377466
rect 199384 377402 199436 377408
rect 199488 377126 199516 377839
rect 199476 377120 199528 377126
rect 199476 377062 199528 377068
rect 199382 371920 199438 371929
rect 199382 371855 199438 371864
rect 198844 354646 198964 354674
rect 198844 353161 198872 354646
rect 198830 353152 198886 353161
rect 198830 353087 198886 353096
rect 198738 291000 198794 291009
rect 198738 290935 198794 290944
rect 198004 271244 198056 271250
rect 198004 271186 198056 271192
rect 197728 270564 197780 270570
rect 197728 270506 197780 270512
rect 197912 270564 197964 270570
rect 197912 270506 197964 270512
rect 197544 253360 197596 253366
rect 197544 253302 197596 253308
rect 197452 165028 197504 165034
rect 197452 164970 197504 164976
rect 197464 57866 197492 164970
rect 197556 146198 197584 253302
rect 197636 253292 197688 253298
rect 197636 253234 197688 253240
rect 197648 146266 197676 253234
rect 197740 165578 197768 270506
rect 198752 183569 198780 290935
rect 198844 246265 198872 353087
rect 199396 296714 199424 371855
rect 199488 370530 199516 377062
rect 199476 370524 199528 370530
rect 199476 370466 199528 370472
rect 199028 296686 199424 296714
rect 198922 291680 198978 291689
rect 198922 291615 198978 291624
rect 198830 246256 198886 246265
rect 198830 246191 198886 246200
rect 198738 183560 198794 183569
rect 198738 183495 198794 183504
rect 198738 182064 198794 182073
rect 198738 181999 198794 182008
rect 197728 165572 197780 165578
rect 197728 165514 197780 165520
rect 197636 146260 197688 146266
rect 197636 146202 197688 146208
rect 197544 146192 197596 146198
rect 197544 146134 197596 146140
rect 198752 74905 198780 181999
rect 198844 139233 198872 246191
rect 198936 184929 198964 291615
rect 199028 288833 199056 296686
rect 199198 292768 199254 292777
rect 199198 292703 199254 292712
rect 199014 288824 199070 288833
rect 199014 288759 199070 288768
rect 198922 184920 198978 184929
rect 198922 184855 198978 184864
rect 198922 183560 198978 183569
rect 198922 183495 198978 183504
rect 198830 139224 198886 139233
rect 198830 139159 198886 139168
rect 198936 76401 198964 183495
rect 199028 182073 199056 288759
rect 199106 288416 199162 288425
rect 199106 288351 199162 288360
rect 199120 287609 199148 288351
rect 199106 287600 199162 287609
rect 199106 287535 199162 287544
rect 199014 182064 199070 182073
rect 199014 181999 199070 182008
rect 199120 180713 199148 287535
rect 199212 209774 199240 292703
rect 199488 291689 199516 370466
rect 199580 369170 199608 400279
rect 199752 398268 199804 398274
rect 199752 398210 199804 398216
rect 199764 394641 199792 398210
rect 199750 394632 199806 394641
rect 199750 394567 199806 394576
rect 199568 369164 199620 369170
rect 199568 369106 199620 369112
rect 199580 364334 199608 369106
rect 199580 364306 199700 364334
rect 199568 362976 199620 362982
rect 199568 362918 199620 362924
rect 199474 291680 199530 291689
rect 199474 291615 199530 291624
rect 199580 288425 199608 362918
rect 199672 292777 199700 364306
rect 199764 363662 199792 394567
rect 200132 380322 200160 484078
rect 200776 480254 200804 488022
rect 201408 485580 201460 485586
rect 201408 485522 201460 485528
rect 200224 480226 200804 480254
rect 200120 380316 200172 380322
rect 200120 380258 200172 380264
rect 200224 380254 200252 480226
rect 200948 475652 201000 475658
rect 200948 475594 201000 475600
rect 200396 471504 200448 471510
rect 200396 471446 200448 471452
rect 200304 465996 200356 466002
rect 200304 465938 200356 465944
rect 200212 380248 200264 380254
rect 200212 380190 200264 380196
rect 199844 378140 199896 378146
rect 199844 378082 199896 378088
rect 199752 363656 199804 363662
rect 199752 363598 199804 363604
rect 199764 362982 199792 363598
rect 199752 362976 199804 362982
rect 199752 362918 199804 362924
rect 199856 362250 199884 378082
rect 199764 362234 199884 362250
rect 199752 362228 199884 362234
rect 199804 362222 199884 362228
rect 199752 362170 199804 362176
rect 199658 292768 199714 292777
rect 199658 292703 199714 292712
rect 199764 291009 199792 362170
rect 200120 358080 200172 358086
rect 200120 358022 200172 358028
rect 199750 291000 199806 291009
rect 199750 290935 199806 290944
rect 199566 288416 199622 288425
rect 199566 288351 199622 288360
rect 200132 271318 200160 358022
rect 200316 271386 200344 465938
rect 200408 377262 200436 471446
rect 200488 471436 200540 471442
rect 200488 471378 200540 471384
rect 200396 377256 200448 377262
rect 200396 377198 200448 377204
rect 200500 377194 200528 471378
rect 200856 468308 200908 468314
rect 200856 468250 200908 468256
rect 200764 467492 200816 467498
rect 200764 467434 200816 467440
rect 200580 465044 200632 465050
rect 200580 464986 200632 464992
rect 200592 380458 200620 464986
rect 200776 389162 200804 467434
rect 200764 389156 200816 389162
rect 200764 389098 200816 389104
rect 200580 380452 200632 380458
rect 200580 380394 200632 380400
rect 200488 377188 200540 377194
rect 200488 377130 200540 377136
rect 200764 359508 200816 359514
rect 200764 359450 200816 359456
rect 200776 282198 200804 359450
rect 200764 282192 200816 282198
rect 200764 282134 200816 282140
rect 200304 271380 200356 271386
rect 200304 271322 200356 271328
rect 200120 271312 200172 271318
rect 200120 271254 200172 271260
rect 200776 253230 200804 282134
rect 200868 272542 200896 468250
rect 200960 284306 200988 475594
rect 201420 379234 201448 485522
rect 201500 484968 201552 484974
rect 201498 484936 201500 484945
rect 201552 484936 201554 484945
rect 201498 484871 201554 484880
rect 201500 483540 201552 483546
rect 201500 483482 201552 483488
rect 201408 379228 201460 379234
rect 201408 379170 201460 379176
rect 201420 378894 201448 379170
rect 201408 378888 201460 378894
rect 201408 378830 201460 378836
rect 201512 378146 201540 483482
rect 201604 380186 201632 488022
rect 201696 488022 201986 488050
rect 202462 488022 202736 488050
rect 202922 488022 203012 488050
rect 203290 488022 203656 488050
rect 201696 483546 201724 488022
rect 202236 485172 202288 485178
rect 202236 485114 202288 485120
rect 201684 483540 201736 483546
rect 201684 483482 201736 483488
rect 201776 482452 201828 482458
rect 201776 482394 201828 482400
rect 201684 468512 201736 468518
rect 201684 468454 201736 468460
rect 201592 380180 201644 380186
rect 201592 380122 201644 380128
rect 201500 378140 201552 378146
rect 201500 378082 201552 378088
rect 201408 360256 201460 360262
rect 201408 360198 201460 360204
rect 201420 359514 201448 360198
rect 201408 359508 201460 359514
rect 201408 359450 201460 359456
rect 200948 284300 201000 284306
rect 200948 284242 201000 284248
rect 200856 272536 200908 272542
rect 200856 272478 200908 272484
rect 201696 271862 201724 468454
rect 201788 376310 201816 482394
rect 202144 474360 202196 474366
rect 202144 474302 202196 474308
rect 201868 471096 201920 471102
rect 201868 471038 201920 471044
rect 201880 380050 201908 471038
rect 201868 380044 201920 380050
rect 201868 379986 201920 379992
rect 201776 376304 201828 376310
rect 201776 376246 201828 376252
rect 201684 271856 201736 271862
rect 201684 271798 201736 271804
rect 202156 271726 202184 474302
rect 202144 271720 202196 271726
rect 202144 271662 202196 271668
rect 200764 253224 200816 253230
rect 200764 253166 200816 253172
rect 199212 209746 199332 209774
rect 199304 186425 199332 209746
rect 199290 186416 199346 186425
rect 199290 186351 199346 186360
rect 199198 184920 199254 184929
rect 199198 184855 199254 184864
rect 199106 180704 199162 180713
rect 199106 180639 199162 180648
rect 199120 161474 199148 180639
rect 199028 161446 199148 161474
rect 198922 76392 198978 76401
rect 198922 76327 198978 76336
rect 198738 74896 198794 74905
rect 198738 74831 198794 74840
rect 199028 73681 199056 161446
rect 199212 77761 199240 184855
rect 199304 79393 199332 186351
rect 200776 175234 200804 253166
rect 200764 175228 200816 175234
rect 200764 175170 200816 175176
rect 201500 175228 201552 175234
rect 201500 175170 201552 175176
rect 201512 145586 201540 175170
rect 202248 166462 202276 485114
rect 202708 485042 202736 488022
rect 202696 485036 202748 485042
rect 202696 484978 202748 484984
rect 202880 471300 202932 471306
rect 202880 471242 202932 471248
rect 202328 469872 202380 469878
rect 202328 469814 202380 469820
rect 202236 166456 202288 166462
rect 202236 166398 202288 166404
rect 202340 164966 202368 469814
rect 202512 467424 202564 467430
rect 202512 467366 202564 467372
rect 202420 466404 202472 466410
rect 202420 466346 202472 466352
rect 202432 272882 202460 466346
rect 202524 376174 202552 467366
rect 202786 379536 202842 379545
rect 202786 379471 202842 379480
rect 202696 379432 202748 379438
rect 202696 379374 202748 379380
rect 202708 378486 202736 379374
rect 202696 378480 202748 378486
rect 202696 378422 202748 378428
rect 202512 376168 202564 376174
rect 202512 376110 202564 376116
rect 202420 272876 202472 272882
rect 202420 272818 202472 272824
rect 202708 268394 202736 378422
rect 202696 268388 202748 268394
rect 202696 268330 202748 268336
rect 202328 164960 202380 164966
rect 202328 164902 202380 164908
rect 201500 145580 201552 145586
rect 201500 145522 201552 145528
rect 199290 79384 199346 79393
rect 199290 79319 199346 79328
rect 199198 77752 199254 77761
rect 199198 77687 199254 77696
rect 199014 73672 199070 73681
rect 199014 73607 199070 73616
rect 202800 58886 202828 379471
rect 202892 271658 202920 471242
rect 202984 380458 203012 488022
rect 203628 486538 203656 488022
rect 203616 486532 203668 486538
rect 203616 486474 203668 486480
rect 203720 484362 203748 488036
rect 203812 488022 204194 488050
rect 204364 488022 204654 488050
rect 204732 488022 205022 488050
rect 205192 488022 205482 488050
rect 205958 488022 206048 488050
rect 203708 484356 203760 484362
rect 203708 484298 203760 484304
rect 203812 484208 203840 488022
rect 204260 486668 204312 486674
rect 204260 486610 204312 486616
rect 204272 485602 204300 486610
rect 204180 485574 204300 485602
rect 204180 485330 204208 485574
rect 204180 485302 204300 485330
rect 203076 484180 203840 484208
rect 202972 380452 203024 380458
rect 202972 380394 203024 380400
rect 203076 380361 203104 484180
rect 203616 482792 203668 482798
rect 203616 482734 203668 482740
rect 203156 482384 203208 482390
rect 203156 482326 203208 482332
rect 203168 380526 203196 482326
rect 203524 478236 203576 478242
rect 203524 478178 203576 478184
rect 203248 465860 203300 465866
rect 203248 465802 203300 465808
rect 203156 380520 203208 380526
rect 203156 380462 203208 380468
rect 203062 380352 203118 380361
rect 203062 380287 203118 380296
rect 203260 380118 203288 465802
rect 203248 380112 203300 380118
rect 203248 380054 203300 380060
rect 202880 271652 202932 271658
rect 202880 271594 202932 271600
rect 203536 164898 203564 478178
rect 203628 271386 203656 482734
rect 203708 471232 203760 471238
rect 203708 471174 203760 471180
rect 203720 272814 203748 471174
rect 203800 466132 203852 466138
rect 203800 466074 203852 466080
rect 203812 282878 203840 466074
rect 203892 465520 203944 465526
rect 203892 465462 203944 465468
rect 203904 376582 203932 465462
rect 203892 376576 203944 376582
rect 203892 376518 203944 376524
rect 203800 282872 203852 282878
rect 203800 282814 203852 282820
rect 203708 272808 203760 272814
rect 203708 272750 203760 272756
rect 204272 271590 204300 485302
rect 204364 380633 204392 488022
rect 204444 485444 204496 485450
rect 204444 485386 204496 485392
rect 204456 485217 204484 485386
rect 204442 485208 204498 485217
rect 204442 485143 204498 485152
rect 204444 484152 204496 484158
rect 204732 484106 204760 488022
rect 205192 484158 205220 488022
rect 205824 487076 205876 487082
rect 205824 487018 205876 487024
rect 205640 486600 205692 486606
rect 205640 486542 205692 486548
rect 205456 485172 205508 485178
rect 205456 485114 205508 485120
rect 204444 484094 204496 484100
rect 204456 411942 204484 484094
rect 204548 484078 204760 484106
rect 205180 484152 205232 484158
rect 205180 484094 205232 484100
rect 204548 477018 204576 484078
rect 205180 483812 205232 483818
rect 205180 483754 205232 483760
rect 204628 482316 204680 482322
rect 204628 482258 204680 482264
rect 204536 477012 204588 477018
rect 204536 476954 204588 476960
rect 204444 411936 204496 411942
rect 204444 411878 204496 411884
rect 204350 380624 204406 380633
rect 204350 380559 204406 380568
rect 204364 380526 204392 380559
rect 204352 380520 204404 380526
rect 204352 380462 204404 380468
rect 204640 380390 204668 482258
rect 204902 471336 204958 471345
rect 204902 471271 204958 471280
rect 204628 380384 204680 380390
rect 204628 380326 204680 380332
rect 204260 271584 204312 271590
rect 204260 271526 204312 271532
rect 203616 271380 203668 271386
rect 203616 271322 203668 271328
rect 204916 166666 204944 471271
rect 205088 469940 205140 469946
rect 205088 469882 205140 469888
rect 204994 466168 205050 466177
rect 204994 466103 205050 466112
rect 204904 166660 204956 166666
rect 204904 166602 204956 166608
rect 205008 166598 205036 466103
rect 205100 178022 205128 469882
rect 205192 271522 205220 483754
rect 205272 464704 205324 464710
rect 205272 464646 205324 464652
rect 205284 272678 205312 464646
rect 205468 378826 205496 485114
rect 205546 411360 205602 411369
rect 205546 411295 205602 411304
rect 205456 378820 205508 378826
rect 205456 378762 205508 378768
rect 205272 272672 205324 272678
rect 205272 272614 205324 272620
rect 205180 271516 205232 271522
rect 205180 271458 205232 271464
rect 205088 178016 205140 178022
rect 205088 177958 205140 177964
rect 204996 166592 205048 166598
rect 204996 166534 205048 166540
rect 203524 164892 203576 164898
rect 203524 164834 203576 164840
rect 204904 145580 204956 145586
rect 204904 145522 204956 145528
rect 204916 67658 204944 145522
rect 204904 67652 204956 67658
rect 204904 67594 204956 67600
rect 202788 58880 202840 58886
rect 202788 58822 202840 58828
rect 204916 57934 204944 67594
rect 205560 59090 205588 411295
rect 205652 271794 205680 486542
rect 205836 480978 205864 487018
rect 206020 485774 206048 488022
rect 206112 488022 206402 488050
rect 206480 488022 206862 488050
rect 207246 488022 207520 488050
rect 206112 487082 206140 488022
rect 206100 487076 206152 487082
rect 206100 487018 206152 487024
rect 206020 485746 206140 485774
rect 205744 480950 205864 480978
rect 205744 413302 205772 480950
rect 205824 480888 205876 480894
rect 205824 480830 205876 480836
rect 205836 416770 205864 480830
rect 206112 475386 206140 485746
rect 206192 485512 206244 485518
rect 206192 485454 206244 485460
rect 206204 485217 206232 485454
rect 206190 485208 206246 485217
rect 206190 485143 206246 485152
rect 206480 480894 206508 488022
rect 206468 480888 206520 480894
rect 206468 480830 206520 480836
rect 207204 480888 207256 480894
rect 207204 480830 207256 480836
rect 207112 477420 207164 477426
rect 207112 477362 207164 477368
rect 206376 475516 206428 475522
rect 206376 475458 206428 475464
rect 206100 475380 206152 475386
rect 206100 475322 206152 475328
rect 205916 471164 205968 471170
rect 205916 471106 205968 471112
rect 205824 416764 205876 416770
rect 205824 416706 205876 416712
rect 205732 413296 205784 413302
rect 205732 413238 205784 413244
rect 205732 411936 205784 411942
rect 205732 411878 205784 411884
rect 205744 410582 205772 411878
rect 205732 410576 205784 410582
rect 205732 410518 205784 410524
rect 205928 380934 205956 471106
rect 206284 389224 206336 389230
rect 206284 389166 206336 389172
rect 206190 381032 206246 381041
rect 206190 380967 206246 380976
rect 205916 380928 205968 380934
rect 205916 380870 205968 380876
rect 205640 271788 205692 271794
rect 205640 271730 205692 271736
rect 205548 59084 205600 59090
rect 205548 59026 205600 59032
rect 204904 57928 204956 57934
rect 204904 57870 204956 57876
rect 206204 57866 206232 380967
rect 206296 360262 206324 389166
rect 206284 360256 206336 360262
rect 206284 360198 206336 360204
rect 206388 165170 206416 475458
rect 206560 471980 206612 471986
rect 206560 471922 206612 471928
rect 206466 466032 206522 466041
rect 206466 465967 206522 465976
rect 206480 166530 206508 465967
rect 206572 272610 206600 471922
rect 206652 469056 206704 469062
rect 206652 468998 206704 469004
rect 206560 272604 206612 272610
rect 206560 272546 206612 272552
rect 206664 271182 206692 468998
rect 207020 466472 207072 466478
rect 207020 466414 207072 466420
rect 206744 466200 206796 466206
rect 206744 466142 206796 466148
rect 206756 273290 206784 466142
rect 206836 417444 206888 417450
rect 206836 417386 206888 417392
rect 206848 378593 206876 417386
rect 206928 414724 206980 414730
rect 206928 414666 206980 414672
rect 206940 379438 206968 414666
rect 207032 390522 207060 466414
rect 207020 390516 207072 390522
rect 207020 390458 207072 390464
rect 207032 389230 207060 390458
rect 207020 389224 207072 389230
rect 207020 389166 207072 389172
rect 207124 379914 207152 477362
rect 207216 417518 207244 480830
rect 207296 474088 207348 474094
rect 207296 474030 207348 474036
rect 207204 417512 207256 417518
rect 207204 417454 207256 417460
rect 207308 380594 207336 474030
rect 207388 465792 207440 465798
rect 207388 465734 207440 465740
rect 207400 380662 207428 465734
rect 207492 465050 207520 488022
rect 207584 488022 207690 488050
rect 207768 488022 208150 488050
rect 208626 488022 208992 488050
rect 207584 480894 207612 488022
rect 207572 480888 207624 480894
rect 207572 480830 207624 480836
rect 207664 479596 207716 479602
rect 207664 479538 207716 479544
rect 207480 465044 207532 465050
rect 207480 464986 207532 464992
rect 207388 380656 207440 380662
rect 207388 380598 207440 380604
rect 207296 380588 207348 380594
rect 207296 380530 207348 380536
rect 207112 379908 207164 379914
rect 207112 379850 207164 379856
rect 206928 379432 206980 379438
rect 206928 379374 206980 379380
rect 206834 378584 206890 378593
rect 206834 378519 206890 378528
rect 207124 376650 207152 379850
rect 207570 379128 207626 379137
rect 207570 379063 207626 379072
rect 207112 376644 207164 376650
rect 207112 376586 207164 376592
rect 206744 273284 206796 273290
rect 206744 273226 206796 273232
rect 206652 271176 206704 271182
rect 206652 271118 206704 271124
rect 207584 270337 207612 379063
rect 207570 270328 207626 270337
rect 207570 270263 207626 270272
rect 207676 175234 207704 479538
rect 207768 477426 207796 488022
rect 208308 485444 208360 485450
rect 208308 485386 208360 485392
rect 207756 477420 207808 477426
rect 207756 477362 207808 477368
rect 207756 476944 207808 476950
rect 207756 476886 207808 476892
rect 207768 271017 207796 476886
rect 207940 465044 207992 465050
rect 207940 464986 207992 464992
rect 207848 464636 207900 464642
rect 207848 464578 207900 464584
rect 207860 272746 207888 464578
rect 207952 464302 207980 464986
rect 207940 464296 207992 464302
rect 207940 464238 207992 464244
rect 207952 422958 207980 464238
rect 207940 422952 207992 422958
rect 207940 422894 207992 422900
rect 207940 416764 207992 416770
rect 207940 416706 207992 416712
rect 207952 414866 207980 416706
rect 207940 414860 207992 414866
rect 207940 414802 207992 414808
rect 208124 414792 208176 414798
rect 208124 414734 208176 414740
rect 208136 383654 208164 414734
rect 208044 383626 208164 383654
rect 207938 379128 207994 379137
rect 207938 379063 207994 379072
rect 207952 378865 207980 379063
rect 207938 378856 207994 378865
rect 207938 378791 207994 378800
rect 208044 375290 208072 383626
rect 208122 380216 208178 380225
rect 208122 380151 208178 380160
rect 208136 379642 208164 380151
rect 208124 379636 208176 379642
rect 208124 379578 208176 379584
rect 208032 375284 208084 375290
rect 208032 375226 208084 375232
rect 208044 374678 208072 375226
rect 208136 375086 208164 379578
rect 208320 379514 208348 485386
rect 208964 485382 208992 488022
rect 208952 485376 209004 485382
rect 208952 485318 209004 485324
rect 208400 485104 208452 485110
rect 208398 485072 208400 485081
rect 208452 485072 208454 485081
rect 208398 485007 208454 485016
rect 209056 484974 209084 488036
rect 209148 488022 209438 488050
rect 209044 484968 209096 484974
rect 209044 484910 209096 484916
rect 208400 484832 208452 484838
rect 208398 484800 208400 484809
rect 208452 484800 208454 484809
rect 208398 484735 208454 484744
rect 209148 476114 209176 488022
rect 209504 485104 209556 485110
rect 209504 485046 209556 485052
rect 209228 481092 209280 481098
rect 209228 481034 209280 481040
rect 208964 476086 209176 476114
rect 208768 464772 208820 464778
rect 208768 464714 208820 464720
rect 208674 390688 208730 390697
rect 208674 390623 208730 390632
rect 208228 379486 208348 379514
rect 208228 378808 208256 379486
rect 208228 378780 208348 378808
rect 208214 378720 208270 378729
rect 208214 378655 208270 378664
rect 208124 375080 208176 375086
rect 208124 375022 208176 375028
rect 208032 374672 208084 374678
rect 208032 374614 208084 374620
rect 207848 272740 207900 272746
rect 207848 272682 207900 272688
rect 207754 271008 207810 271017
rect 207754 270943 207810 270952
rect 208228 269754 208256 378655
rect 208320 375358 208348 378780
rect 208308 375352 208360 375358
rect 208308 375294 208360 375300
rect 208306 270328 208362 270337
rect 208306 270263 208362 270272
rect 208216 269748 208268 269754
rect 208216 269690 208268 269696
rect 207664 175228 207716 175234
rect 207664 175170 207716 175176
rect 206468 166524 206520 166530
rect 206468 166466 206520 166472
rect 206376 165164 206428 165170
rect 206376 165106 206428 165112
rect 208320 147490 208348 270263
rect 208308 147484 208360 147490
rect 208308 147426 208360 147432
rect 197452 57860 197504 57866
rect 197452 57802 197504 57808
rect 206192 57860 206244 57866
rect 206192 57802 206244 57808
rect 183468 57792 183520 57798
rect 183466 57760 183468 57769
rect 197360 57792 197412 57798
rect 183520 57760 183522 57769
rect 197360 57734 197412 57740
rect 183466 57695 183522 57704
rect 208688 57662 208716 390623
rect 208780 375970 208808 464714
rect 208858 378992 208914 379001
rect 208964 378962 208992 476086
rect 209044 474224 209096 474230
rect 209044 474166 209096 474172
rect 208858 378927 208914 378936
rect 208952 378956 209004 378962
rect 208768 375964 208820 375970
rect 208768 375906 208820 375912
rect 208872 269793 208900 378927
rect 208952 378898 209004 378904
rect 208964 378690 208992 378898
rect 208952 378684 209004 378690
rect 208952 378626 209004 378632
rect 208952 377528 209004 377534
rect 208952 377470 209004 377476
rect 208858 269784 208914 269793
rect 208858 269719 208914 269728
rect 208964 269074 208992 377470
rect 208952 269068 209004 269074
rect 208952 269010 209004 269016
rect 209056 70378 209084 474166
rect 209136 468852 209188 468858
rect 209136 468794 209188 468800
rect 209148 166394 209176 468794
rect 209240 271114 209268 481034
rect 209320 471776 209372 471782
rect 209320 471718 209372 471724
rect 209332 273086 209360 471718
rect 209412 466064 209464 466070
rect 209412 466006 209464 466012
rect 209320 273080 209372 273086
rect 209320 273022 209372 273028
rect 209424 271250 209452 466006
rect 209516 379642 209544 485046
rect 209596 484356 209648 484362
rect 209596 484298 209648 484304
rect 209608 391950 209636 484298
rect 209780 480888 209832 480894
rect 209780 480830 209832 480836
rect 209688 465724 209740 465730
rect 209688 465666 209740 465672
rect 209596 391944 209648 391950
rect 209596 391886 209648 391892
rect 209504 379636 209556 379642
rect 209504 379578 209556 379584
rect 209594 379536 209650 379545
rect 209594 379471 209650 379480
rect 209502 375456 209558 375465
rect 209502 375391 209558 375400
rect 209412 271244 209464 271250
rect 209412 271186 209464 271192
rect 209228 271108 209280 271114
rect 209228 271050 209280 271056
rect 209412 269748 209464 269754
rect 209412 269690 209464 269696
rect 209136 166388 209188 166394
rect 209136 166330 209188 166336
rect 209424 144838 209452 269690
rect 209412 144832 209464 144838
rect 209412 144774 209464 144780
rect 209044 70372 209096 70378
rect 209044 70314 209096 70320
rect 209516 58750 209544 375391
rect 209608 58818 209636 379471
rect 209700 379030 209728 465666
rect 209792 379370 209820 480830
rect 209884 379506 209912 488036
rect 209976 488022 210358 488050
rect 210528 488022 210818 488050
rect 211202 488022 211292 488050
rect 209976 480894 210004 488022
rect 210528 485774 210556 488022
rect 210068 485746 210556 485774
rect 211160 485784 211212 485790
rect 211158 485752 211160 485761
rect 211212 485752 211214 485761
rect 209964 480888 210016 480894
rect 209964 480830 210016 480836
rect 210068 470594 210096 485746
rect 211158 485687 211214 485696
rect 211160 485648 211212 485654
rect 211160 485590 211212 485596
rect 210148 485036 210200 485042
rect 210148 484978 210200 484984
rect 209976 470566 210096 470594
rect 209976 469169 210004 470566
rect 209962 469160 210018 469169
rect 209962 469095 210018 469104
rect 210056 468376 210108 468382
rect 210056 468318 210108 468324
rect 209872 379500 209924 379506
rect 209872 379442 209924 379448
rect 209780 379364 209832 379370
rect 209780 379306 209832 379312
rect 209884 379234 209912 379442
rect 209872 379228 209924 379234
rect 209872 379170 209924 379176
rect 209688 379024 209740 379030
rect 209688 378966 209740 378972
rect 210068 376446 210096 468318
rect 210160 376650 210188 484978
rect 211172 484673 211200 485590
rect 211158 484664 211214 484673
rect 211158 484599 211214 484608
rect 210700 478304 210752 478310
rect 210700 478246 210752 478252
rect 210516 474292 210568 474298
rect 210516 474234 210568 474240
rect 210424 467152 210476 467158
rect 210424 467094 210476 467100
rect 210332 378820 210384 378826
rect 210332 378762 210384 378768
rect 210240 378480 210292 378486
rect 210240 378422 210292 378428
rect 210252 378282 210280 378422
rect 210344 378282 210372 378762
rect 210240 378276 210292 378282
rect 210240 378218 210292 378224
rect 210332 378276 210384 378282
rect 210332 378218 210384 378224
rect 210148 376644 210200 376650
rect 210148 376586 210200 376592
rect 210056 376440 210108 376446
rect 210056 376382 210108 376388
rect 210252 270094 210280 378218
rect 210344 270162 210372 378218
rect 210332 270156 210384 270162
rect 210332 270098 210384 270104
rect 210240 270088 210292 270094
rect 210240 270030 210292 270036
rect 209596 58812 209648 58818
rect 209596 58754 209648 58760
rect 209504 58744 209556 58750
rect 209504 58686 209556 58692
rect 208676 57656 208728 57662
rect 155958 57624 156014 57633
rect 155958 57559 156014 57568
rect 160098 57624 160154 57633
rect 160098 57559 160154 57568
rect 165618 57624 165674 57633
rect 208676 57598 208728 57604
rect 165618 57559 165674 57568
rect 153290 56264 153346 56273
rect 153290 56199 153346 56208
rect 155972 54913 156000 57559
rect 160112 55049 160140 57559
rect 165632 55185 165660 57559
rect 210436 57458 210464 467094
rect 210528 165510 210556 474234
rect 210608 471572 210660 471578
rect 210608 471514 210660 471520
rect 210620 166734 210648 471514
rect 210712 271318 210740 478246
rect 210792 472728 210844 472734
rect 210792 472670 210844 472676
rect 210700 271312 210752 271318
rect 210700 271254 210752 271260
rect 210804 271046 210832 472670
rect 210884 471708 210936 471714
rect 210884 471650 210936 471656
rect 210896 272950 210924 471650
rect 211264 379302 211292 488022
rect 211632 485586 211660 488036
rect 211724 488022 212106 488050
rect 212582 488022 212764 488050
rect 211620 485580 211672 485586
rect 211620 485522 211672 485528
rect 211724 470594 211752 488022
rect 212540 485716 212592 485722
rect 212540 485658 212592 485664
rect 212552 485625 212580 485658
rect 212538 485616 212594 485625
rect 212538 485551 212594 485560
rect 212736 481098 212764 488022
rect 212828 488022 213026 488050
rect 212724 481092 212776 481098
rect 212724 481034 212776 481040
rect 211804 481024 211856 481030
rect 211804 480966 211856 480972
rect 211356 470566 211752 470594
rect 211356 379506 211384 470566
rect 211620 468444 211672 468450
rect 211620 468386 211672 468392
rect 211528 466336 211580 466342
rect 211528 466278 211580 466284
rect 211344 379500 211396 379506
rect 211344 379442 211396 379448
rect 211252 379296 211304 379302
rect 211252 379238 211304 379244
rect 211264 379098 211292 379238
rect 211252 379092 211304 379098
rect 211252 379034 211304 379040
rect 211356 378486 211384 379442
rect 211344 378480 211396 378486
rect 211344 378422 211396 378428
rect 210974 375592 211030 375601
rect 210974 375527 211030 375536
rect 210884 272944 210936 272950
rect 210884 272886 210936 272892
rect 210792 271040 210844 271046
rect 210792 270982 210844 270988
rect 210882 270192 210938 270201
rect 210882 270127 210938 270136
rect 210608 166728 210660 166734
rect 210608 166670 210660 166676
rect 210516 165504 210568 165510
rect 210516 165446 210568 165452
rect 210896 147626 210924 270127
rect 210884 147620 210936 147626
rect 210884 147562 210936 147568
rect 210988 57526 211016 375527
rect 211066 375456 211122 375465
rect 211066 375391 211122 375400
rect 211080 57934 211108 375391
rect 211540 270473 211568 466278
rect 211632 376514 211660 468386
rect 211710 379128 211766 379137
rect 211710 379063 211766 379072
rect 211620 376508 211672 376514
rect 211620 376450 211672 376456
rect 211724 273494 211752 379063
rect 211712 273488 211764 273494
rect 211712 273430 211764 273436
rect 211526 270464 211582 270473
rect 211526 270399 211582 270408
rect 211816 164762 211844 480966
rect 212540 480888 212592 480894
rect 212540 480830 212592 480836
rect 211896 476808 211948 476814
rect 211896 476750 211948 476756
rect 211908 165306 211936 476750
rect 212080 474020 212132 474026
rect 212080 473962 212132 473968
rect 211986 468752 212042 468761
rect 211986 468687 212042 468696
rect 212000 166326 212028 468687
rect 212092 271697 212120 473962
rect 212356 468988 212408 468994
rect 212356 468930 212408 468936
rect 212172 467356 212224 467362
rect 212172 467298 212224 467304
rect 212184 271794 212212 467298
rect 212264 274780 212316 274786
rect 212264 274722 212316 274728
rect 212172 271788 212224 271794
rect 212172 271730 212224 271736
rect 212078 271688 212134 271697
rect 212078 271623 212134 271632
rect 212172 268388 212224 268394
rect 212172 268330 212224 268336
rect 212184 166802 212212 268330
rect 212172 166796 212224 166802
rect 212172 166738 212224 166744
rect 211988 166320 212040 166326
rect 211988 166262 212040 166268
rect 211896 165300 211948 165306
rect 211896 165242 211948 165248
rect 211804 164756 211856 164762
rect 211804 164698 211856 164704
rect 212276 163946 212304 274722
rect 212368 273154 212396 468930
rect 212552 379574 212580 480830
rect 212828 478156 212856 488022
rect 213380 484430 213408 488036
rect 213472 488022 213854 488050
rect 214024 488022 214314 488050
rect 213368 484424 213420 484430
rect 213368 484366 213420 484372
rect 212908 481092 212960 481098
rect 212908 481034 212960 481040
rect 212644 478128 212856 478156
rect 212644 379778 212672 478128
rect 212920 473354 212948 481034
rect 213472 480894 213500 488022
rect 213460 480888 213512 480894
rect 213460 480830 213512 480836
rect 213276 476876 213328 476882
rect 213276 476818 213328 476824
rect 213184 475448 213236 475454
rect 213184 475390 213236 475396
rect 212736 473326 212948 473354
rect 212632 379772 212684 379778
rect 212632 379714 212684 379720
rect 212736 379710 212764 473326
rect 213092 469192 213144 469198
rect 213092 469134 213144 469140
rect 212816 466472 212868 466478
rect 212816 466414 212868 466420
rect 212828 381070 212856 466414
rect 213000 465656 213052 465662
rect 213000 465598 213052 465604
rect 212816 381064 212868 381070
rect 212816 381006 212868 381012
rect 212814 380352 212870 380361
rect 212814 380287 212870 380296
rect 212724 379704 212776 379710
rect 212724 379646 212776 379652
rect 212540 379568 212592 379574
rect 212540 379510 212592 379516
rect 212552 379302 212580 379510
rect 212540 379296 212592 379302
rect 212540 379238 212592 379244
rect 212540 378820 212592 378826
rect 212540 378762 212592 378768
rect 212552 378214 212580 378762
rect 212630 378584 212686 378593
rect 212630 378519 212686 378528
rect 212540 378208 212592 378214
rect 212446 378176 212502 378185
rect 212644 378185 212672 378519
rect 212540 378150 212592 378156
rect 212630 378176 212686 378185
rect 212446 378111 212502 378120
rect 212630 378111 212686 378120
rect 212356 273148 212408 273154
rect 212356 273090 212408 273096
rect 212354 269784 212410 269793
rect 212354 269719 212410 269728
rect 212264 163940 212316 163946
rect 212264 163882 212316 163888
rect 212368 147558 212396 269719
rect 212356 147552 212408 147558
rect 212356 147494 212408 147500
rect 212460 58954 212488 378111
rect 212632 376440 212684 376446
rect 212630 376408 212632 376417
rect 212684 376408 212686 376417
rect 212540 376372 212592 376378
rect 212630 376343 212686 376352
rect 212540 376314 212592 376320
rect 212552 375630 212580 376314
rect 212736 376242 212764 379646
rect 212724 376236 212776 376242
rect 212724 376178 212776 376184
rect 212540 375624 212592 375630
rect 212540 375566 212592 375572
rect 212828 271833 212856 380287
rect 212908 379296 212960 379302
rect 212908 379238 212960 379244
rect 212920 377534 212948 379238
rect 212908 377528 212960 377534
rect 212908 377470 212960 377476
rect 213012 376718 213040 465598
rect 213000 376712 213052 376718
rect 213000 376654 213052 376660
rect 213104 376378 213132 469134
rect 213092 376372 213144 376378
rect 213092 376314 213144 376320
rect 213092 273352 213144 273358
rect 213092 273294 213144 273300
rect 212814 271824 212870 271833
rect 212814 271759 212870 271768
rect 213000 270496 213052 270502
rect 213000 270438 213052 270444
rect 213012 144770 213040 270438
rect 213104 148442 213132 273294
rect 213196 165442 213224 475390
rect 213288 270910 213316 476818
rect 213828 466404 213880 466410
rect 213828 466346 213880 466352
rect 213644 380520 213696 380526
rect 213644 380462 213696 380468
rect 213656 379846 213684 380462
rect 213734 380352 213790 380361
rect 213734 380287 213790 380296
rect 213748 379982 213776 380287
rect 213736 379976 213788 379982
rect 213736 379918 213788 379924
rect 213644 379840 213696 379846
rect 213644 379782 213696 379788
rect 213368 379500 213420 379506
rect 213368 379442 213420 379448
rect 213380 379302 213408 379442
rect 213368 379296 213420 379302
rect 213368 379238 213420 379244
rect 213460 378820 213512 378826
rect 213460 378762 213512 378768
rect 213368 378344 213420 378350
rect 213368 378286 213420 378292
rect 213380 273358 213408 378286
rect 213368 273352 213420 273358
rect 213368 273294 213420 273300
rect 213366 271824 213422 271833
rect 213366 271759 213422 271768
rect 213380 271425 213408 271759
rect 213366 271416 213422 271425
rect 213366 271351 213422 271360
rect 213276 270904 213328 270910
rect 213276 270846 213328 270852
rect 213184 165436 213236 165442
rect 213184 165378 213236 165384
rect 213380 164082 213408 271351
rect 213472 270502 213500 378762
rect 213552 376440 213604 376446
rect 213550 376408 213552 376417
rect 213604 376408 213606 376417
rect 213550 376343 213606 376352
rect 213552 375420 213604 375426
rect 213552 375362 213604 375368
rect 213460 270496 213512 270502
rect 213460 270438 213512 270444
rect 213472 270298 213500 270438
rect 213460 270292 213512 270298
rect 213460 270234 213512 270240
rect 213460 270156 213512 270162
rect 213460 270098 213512 270104
rect 213472 269822 213500 270098
rect 213460 269816 213512 269822
rect 213460 269758 213512 269764
rect 213368 164076 213420 164082
rect 213368 164018 213420 164024
rect 213368 163940 213420 163946
rect 213368 163882 213420 163888
rect 213380 163538 213408 163882
rect 213368 163532 213420 163538
rect 213368 163474 213420 163480
rect 213276 148640 213328 148646
rect 213276 148582 213328 148588
rect 213092 148436 213144 148442
rect 213092 148378 213144 148384
rect 213288 147558 213316 148582
rect 213276 147552 213328 147558
rect 213276 147494 213328 147500
rect 213184 147484 213236 147490
rect 213184 147426 213236 147432
rect 213000 144764 213052 144770
rect 213000 144706 213052 144712
rect 212448 58948 212500 58954
rect 212448 58890 212500 58896
rect 211068 57928 211120 57934
rect 211068 57870 211120 57876
rect 210976 57520 211028 57526
rect 210976 57462 211028 57468
rect 210424 57452 210476 57458
rect 210424 57394 210476 57400
rect 213196 55826 213224 147426
rect 213288 55894 213316 147494
rect 213276 55888 213328 55894
rect 213276 55830 213328 55836
rect 213184 55820 213236 55826
rect 213184 55762 213236 55768
rect 165618 55176 165674 55185
rect 165618 55111 165674 55120
rect 160098 55040 160154 55049
rect 160098 54975 160154 54984
rect 155958 54904 156014 54913
rect 155958 54839 156014 54848
rect 92480 54742 92532 54748
rect 118698 54768 118754 54777
rect 89812 54732 89864 54738
rect 118698 54703 118754 54712
rect 89812 54674 89864 54680
rect 80060 54664 80112 54670
rect 80060 54606 80112 54612
rect 213380 54466 213408 163474
rect 213472 148374 213500 269758
rect 213564 268666 213592 375362
rect 213656 269006 213684 379782
rect 213840 379273 213868 466346
rect 213920 379772 213972 379778
rect 213920 379714 213972 379720
rect 213826 379264 213882 379273
rect 213826 379199 213882 379208
rect 213840 378321 213868 379199
rect 213826 378312 213882 378321
rect 213826 378247 213882 378256
rect 213932 377482 213960 379714
rect 213840 377454 213960 377482
rect 213840 377346 213868 377454
rect 214024 377346 214052 488022
rect 214760 484537 214788 488036
rect 214852 488022 215234 488050
rect 215312 488022 215602 488050
rect 215680 488022 216062 488050
rect 216232 488022 216522 488050
rect 216876 488022 216982 488050
rect 214746 484528 214802 484537
rect 214746 484463 214802 484472
rect 214852 483800 214880 488022
rect 214932 484424 214984 484430
rect 214932 484366 214984 484372
rect 214208 483772 214880 483800
rect 214208 383654 214236 483772
rect 214564 483676 214616 483682
rect 214564 483618 214616 483624
rect 214208 383626 214512 383654
rect 214104 379500 214156 379506
rect 214104 379442 214156 379448
rect 214116 378418 214144 379442
rect 214104 378412 214156 378418
rect 214104 378354 214156 378360
rect 213748 377318 213868 377346
rect 213932 377318 214052 377346
rect 213748 376038 213776 377318
rect 213826 376816 213882 376825
rect 213826 376751 213882 376760
rect 213736 376032 213788 376038
rect 213736 375974 213788 375980
rect 213748 375426 213776 375974
rect 213736 375420 213788 375426
rect 213736 375362 213788 375368
rect 213736 274712 213788 274718
rect 213736 274654 213788 274660
rect 213748 273358 213776 274654
rect 213736 273352 213788 273358
rect 213736 273294 213788 273300
rect 213644 269000 213696 269006
rect 213644 268942 213696 268948
rect 213552 268660 213604 268666
rect 213552 268602 213604 268608
rect 213748 151814 213776 273294
rect 213564 151786 213776 151814
rect 213564 149054 213592 151786
rect 213552 149048 213604 149054
rect 213552 148990 213604 148996
rect 213460 148368 213512 148374
rect 213460 148310 213512 148316
rect 213458 145616 213514 145625
rect 213458 145551 213514 145560
rect 213472 144838 213500 145551
rect 213460 144832 213512 144838
rect 213460 144774 213512 144780
rect 213368 54460 213420 54466
rect 213368 54402 213420 54408
rect 213472 54398 213500 144774
rect 213564 56506 213592 148990
rect 213736 148504 213788 148510
rect 213736 148446 213788 148452
rect 213748 147490 213776 148446
rect 213736 147484 213788 147490
rect 213736 147426 213788 147432
rect 213736 146328 213788 146334
rect 213736 146270 213788 146276
rect 213552 56500 213604 56506
rect 213552 56442 213604 56448
rect 213748 55185 213776 146270
rect 213840 59022 213868 376751
rect 213932 376514 213960 377318
rect 213920 376508 213972 376514
rect 213920 376450 213972 376456
rect 213932 376106 213960 376450
rect 213920 376100 213972 376106
rect 213920 376042 213972 376048
rect 214116 274718 214144 378354
rect 214380 375624 214432 375630
rect 214380 375566 214432 375572
rect 214104 274712 214156 274718
rect 214104 274654 214156 274660
rect 214196 273488 214248 273494
rect 214196 273430 214248 273436
rect 214208 146305 214236 273430
rect 214288 269272 214340 269278
rect 214288 269214 214340 269220
rect 214194 146296 214250 146305
rect 214194 146231 214250 146240
rect 214300 144906 214328 269214
rect 214392 268802 214420 375566
rect 214484 375154 214512 383626
rect 214472 375148 214524 375154
rect 214472 375090 214524 375096
rect 214380 268796 214432 268802
rect 214380 268738 214432 268744
rect 214484 252550 214512 375090
rect 214472 252544 214524 252550
rect 214472 252486 214524 252492
rect 214576 164694 214604 483618
rect 214656 482656 214708 482662
rect 214656 482598 214708 482604
rect 214668 165374 214696 482598
rect 214748 468920 214800 468926
rect 214748 468862 214800 468868
rect 214760 271658 214788 468862
rect 214840 465928 214892 465934
rect 214840 465870 214892 465876
rect 214748 271652 214800 271658
rect 214748 271594 214800 271600
rect 214852 270978 214880 465870
rect 214944 380050 214972 484366
rect 215024 471912 215076 471918
rect 215024 471854 215076 471860
rect 214932 380044 214984 380050
rect 214932 379986 214984 379992
rect 214944 375630 214972 379986
rect 215036 375902 215064 471854
rect 215024 375896 215076 375902
rect 215024 375838 215076 375844
rect 214932 375624 214984 375630
rect 214932 375566 214984 375572
rect 215114 375592 215170 375601
rect 215114 375527 215170 375536
rect 214932 358216 214984 358222
rect 214932 358158 214984 358164
rect 214840 270972 214892 270978
rect 214840 270914 214892 270920
rect 214944 270201 214972 358158
rect 214930 270192 214986 270201
rect 214930 270127 214986 270136
rect 214840 268864 214892 268870
rect 214840 268806 214892 268812
rect 214748 252544 214800 252550
rect 214748 252486 214800 252492
rect 214760 252414 214788 252486
rect 214748 252408 214800 252414
rect 214748 252350 214800 252356
rect 214656 165368 214708 165374
rect 214656 165310 214708 165316
rect 214564 164688 214616 164694
rect 214564 164630 214616 164636
rect 214760 162790 214788 252350
rect 214748 162784 214800 162790
rect 214748 162726 214800 162732
rect 214656 162444 214708 162450
rect 214656 162386 214708 162392
rect 214564 147620 214616 147626
rect 214564 147562 214616 147568
rect 214472 146192 214524 146198
rect 214472 146134 214524 146140
rect 214288 144900 214340 144906
rect 214288 144842 214340 144848
rect 214484 59634 214512 146134
rect 214472 59628 214524 59634
rect 214472 59570 214524 59576
rect 213828 59016 213880 59022
rect 213828 58958 213880 58964
rect 213734 55176 213790 55185
rect 213734 55111 213790 55120
rect 213460 54392 213512 54398
rect 213460 54334 213512 54340
rect 214576 54330 214604 147562
rect 214668 59226 214696 162386
rect 214656 59220 214708 59226
rect 214656 59162 214708 59168
rect 214760 59158 214788 162726
rect 214852 145654 214880 268806
rect 214932 148572 214984 148578
rect 214932 148514 214984 148520
rect 214944 147626 214972 148514
rect 215024 148436 215076 148442
rect 215024 148378 215076 148384
rect 214932 147620 214984 147626
rect 214932 147562 214984 147568
rect 214930 146296 214986 146305
rect 214930 146231 214986 146240
rect 214840 145648 214892 145654
rect 214840 145590 214892 145596
rect 214748 59152 214800 59158
rect 214748 59094 214800 59100
rect 214852 54602 214880 145590
rect 214944 55049 214972 146231
rect 215036 56370 215064 148378
rect 215128 57730 215156 375527
rect 215206 375456 215262 375465
rect 215206 375391 215262 375400
rect 215116 57724 215168 57730
rect 215116 57666 215168 57672
rect 215220 57322 215248 375391
rect 215312 375222 215340 488022
rect 215392 484152 215444 484158
rect 215392 484094 215444 484100
rect 215404 377942 215432 484094
rect 215680 470594 215708 488022
rect 216232 484158 216260 488022
rect 216220 484152 216272 484158
rect 216220 484094 216272 484100
rect 216772 484152 216824 484158
rect 216772 484094 216824 484100
rect 215944 483744 215996 483750
rect 215944 483686 215996 483692
rect 215496 470566 215708 470594
rect 215496 380905 215524 470566
rect 215852 466268 215904 466274
rect 215852 466210 215904 466216
rect 215482 380896 215538 380905
rect 215482 380831 215538 380840
rect 215392 377936 215444 377942
rect 215392 377878 215444 377884
rect 215760 377936 215812 377942
rect 215760 377878 215812 377884
rect 215772 377534 215800 377878
rect 215760 377528 215812 377534
rect 215760 377470 215812 377476
rect 215864 376106 215892 466210
rect 215852 376100 215904 376106
rect 215852 376042 215904 376048
rect 215300 375216 215352 375222
rect 215300 375158 215352 375164
rect 215852 358692 215904 358698
rect 215852 358634 215904 358640
rect 215760 357604 215812 357610
rect 215760 357546 215812 357552
rect 215772 277394 215800 357546
rect 215680 277366 215800 277394
rect 215680 274786 215708 277366
rect 215668 274780 215720 274786
rect 215668 274722 215720 274728
rect 215680 273970 215708 274722
rect 215668 273964 215720 273970
rect 215668 273906 215720 273912
rect 215666 273320 215722 273329
rect 215666 273255 215722 273264
rect 215680 57594 215708 273255
rect 215864 271930 215892 358634
rect 215852 271924 215904 271930
rect 215852 271866 215904 271872
rect 215852 269000 215904 269006
rect 215852 268942 215904 268948
rect 215864 268734 215892 268942
rect 215852 268728 215904 268734
rect 215852 268670 215904 268676
rect 215760 252476 215812 252482
rect 215760 252418 215812 252424
rect 215772 162450 215800 252418
rect 215760 162444 215812 162450
rect 215760 162386 215812 162392
rect 215864 146198 215892 268670
rect 215956 164830 215984 483686
rect 216036 482724 216088 482730
rect 216036 482666 216088 482672
rect 216048 165578 216076 482666
rect 216220 472660 216272 472666
rect 216220 472602 216272 472608
rect 216126 465896 216182 465905
rect 216126 465831 216182 465840
rect 216036 165572 216088 165578
rect 216036 165514 216088 165520
rect 216140 165034 216168 465831
rect 216232 271590 216260 472602
rect 216312 471640 216364 471646
rect 216312 471582 216364 471588
rect 216324 273018 216352 471582
rect 216678 417888 216734 417897
rect 216678 417823 216734 417832
rect 216692 417518 216720 417823
rect 216680 417512 216732 417518
rect 216680 417454 216732 417460
rect 216692 402974 216720 417454
rect 216784 414730 216812 484094
rect 216876 414798 216904 488022
rect 217428 485450 217456 488036
rect 217520 488022 217810 488050
rect 218286 488022 218376 488050
rect 218746 488022 219112 488050
rect 217416 485444 217468 485450
rect 217416 485386 217468 485392
rect 217416 485308 217468 485314
rect 217416 485250 217468 485256
rect 217428 480254 217456 485250
rect 217520 484158 217548 488022
rect 218152 485376 218204 485382
rect 218152 485318 218204 485324
rect 217508 484152 217560 484158
rect 217508 484094 217560 484100
rect 217428 480226 217548 480254
rect 217324 477012 217376 477018
rect 217324 476954 217376 476960
rect 217140 414860 217192 414866
rect 217140 414802 217192 414808
rect 216864 414792 216916 414798
rect 217152 414769 217180 414802
rect 216864 414734 216916 414740
rect 217138 414760 217194 414769
rect 216772 414724 216824 414730
rect 217138 414695 217194 414704
rect 216772 414666 216824 414672
rect 216862 413808 216918 413817
rect 216862 413743 216918 413752
rect 216876 413302 216904 413743
rect 216864 413296 216916 413302
rect 216864 413238 216916 413244
rect 216770 410952 216826 410961
rect 216770 410887 216826 410896
rect 216784 410582 216812 410887
rect 216772 410576 216824 410582
rect 216772 410518 216824 410524
rect 216692 402946 216812 402974
rect 216680 391944 216732 391950
rect 216680 391886 216732 391892
rect 216692 390969 216720 391886
rect 216678 390960 216734 390969
rect 216678 390895 216734 390904
rect 216680 390516 216732 390522
rect 216680 390458 216732 390464
rect 216692 389337 216720 390458
rect 216678 389328 216734 389337
rect 216678 389263 216734 389272
rect 216680 389156 216732 389162
rect 216680 389098 216732 389104
rect 216692 389065 216720 389098
rect 216678 389056 216734 389065
rect 216678 388991 216734 389000
rect 216586 380896 216642 380905
rect 216586 380831 216642 380840
rect 216496 379908 216548 379914
rect 216496 379850 216548 379856
rect 216404 376508 216456 376514
rect 216404 376450 216456 376456
rect 216416 375630 216444 376450
rect 216404 375624 216456 375630
rect 216404 375566 216456 375572
rect 216312 273012 216364 273018
rect 216312 272954 216364 272960
rect 216312 271924 216364 271930
rect 216312 271866 216364 271872
rect 216220 271584 216272 271590
rect 216220 271526 216272 271532
rect 216220 269000 216272 269006
rect 216220 268942 216272 268948
rect 216128 165028 216180 165034
rect 216128 164970 216180 164976
rect 215944 164824 215996 164830
rect 215944 164766 215996 164772
rect 215944 148368 215996 148374
rect 215944 148310 215996 148316
rect 215852 146192 215904 146198
rect 215852 146134 215904 146140
rect 215760 146056 215812 146062
rect 215760 145998 215812 146004
rect 215668 57588 215720 57594
rect 215668 57530 215720 57536
rect 215208 57316 215260 57322
rect 215208 57258 215260 57264
rect 215024 56364 215076 56370
rect 215024 56306 215076 56312
rect 215772 56166 215800 145998
rect 215760 56160 215812 56166
rect 215760 56102 215812 56108
rect 215956 55146 215984 148310
rect 216128 145852 216180 145858
rect 216128 145794 216180 145800
rect 216036 145036 216088 145042
rect 216036 144978 216088 144984
rect 216048 144770 216076 144978
rect 216036 144764 216088 144770
rect 216036 144706 216088 144712
rect 216048 55962 216076 144706
rect 216140 56030 216168 145794
rect 216232 145722 216260 268942
rect 216324 148986 216352 271866
rect 216416 252482 216444 375566
rect 216508 269006 216536 379850
rect 216600 375698 216628 380831
rect 216678 380760 216734 380769
rect 216678 380695 216734 380704
rect 216692 379681 216720 380695
rect 216678 379672 216734 379681
rect 216678 379607 216734 379616
rect 216588 375692 216640 375698
rect 216588 375634 216640 375640
rect 216588 375216 216640 375222
rect 216588 375158 216640 375164
rect 216600 269686 216628 375158
rect 216692 373994 216720 379607
rect 216784 375834 216812 402946
rect 216876 380866 216904 413238
rect 216956 410576 217008 410582
rect 216956 410518 217008 410524
rect 216864 380860 216916 380866
rect 216864 380802 216916 380808
rect 216876 379488 216904 380802
rect 216968 380730 216996 410518
rect 216956 380724 217008 380730
rect 216956 380666 217008 380672
rect 216968 379642 216996 380666
rect 217152 380089 217180 414695
rect 217230 411360 217286 411369
rect 217230 411295 217286 411304
rect 217244 402974 217272 411295
rect 217336 409193 217364 476954
rect 217416 471844 217468 471850
rect 217416 471786 217468 471792
rect 217322 409184 217378 409193
rect 217322 409119 217378 409128
rect 217244 402946 217364 402974
rect 217336 380798 217364 402946
rect 217428 382294 217456 471786
rect 217416 382288 217468 382294
rect 217416 382230 217468 382236
rect 217324 380792 217376 380798
rect 217324 380734 217376 380740
rect 217138 380080 217194 380089
rect 217138 380015 217194 380024
rect 216956 379636 217008 379642
rect 216956 379578 217008 379584
rect 217152 379545 217180 380015
rect 217138 379536 217194 379545
rect 216876 379460 216996 379488
rect 217138 379471 217194 379480
rect 216772 375828 216824 375834
rect 216772 375770 216824 375776
rect 216968 373994 216996 379460
rect 217232 375692 217284 375698
rect 217232 375634 217284 375640
rect 216692 373966 216904 373994
rect 216968 373966 217088 373994
rect 216876 306374 216904 373966
rect 217060 307737 217088 373966
rect 217138 310040 217194 310049
rect 217138 309975 217194 309984
rect 217046 307728 217102 307737
rect 217046 307663 217102 307672
rect 216876 306346 216996 306374
rect 216770 305008 216826 305017
rect 216770 304943 216826 304952
rect 216680 284300 216732 284306
rect 216680 284242 216732 284248
rect 216692 284073 216720 284242
rect 216678 284064 216734 284073
rect 216678 283999 216734 284008
rect 216678 282296 216734 282305
rect 216678 282231 216734 282240
rect 216692 282198 216720 282231
rect 216680 282192 216732 282198
rect 216680 282134 216732 282140
rect 216588 269680 216640 269686
rect 216588 269622 216640 269628
rect 216496 269000 216548 269006
rect 216496 268942 216548 268948
rect 216404 252476 216456 252482
rect 216404 252418 216456 252424
rect 216404 251864 216456 251870
rect 216404 251806 216456 251812
rect 216416 162722 216444 251806
rect 216404 162716 216456 162722
rect 216404 162658 216456 162664
rect 216312 148980 216364 148986
rect 216312 148922 216364 148928
rect 216220 145716 216272 145722
rect 216220 145658 216272 145664
rect 216324 56438 216352 148922
rect 216416 58614 216444 162658
rect 216600 146033 216628 269622
rect 216784 198121 216812 304943
rect 216968 302161 216996 306346
rect 216954 302152 217010 302161
rect 216954 302087 217010 302096
rect 216864 282872 216916 282878
rect 216864 282814 216916 282820
rect 216876 282169 216904 282814
rect 216862 282160 216918 282169
rect 216862 282095 216918 282104
rect 216864 270428 216916 270434
rect 216864 270370 216916 270376
rect 216770 198112 216826 198121
rect 216770 198047 216826 198056
rect 216770 197024 216826 197033
rect 216770 196959 216826 196968
rect 216680 178016 216732 178022
rect 216680 177958 216732 177964
rect 216692 177041 216720 177958
rect 216678 177032 216734 177041
rect 216678 176967 216734 176976
rect 216678 175400 216734 175409
rect 216678 175335 216734 175344
rect 216692 175302 216720 175335
rect 216680 175296 216732 175302
rect 216680 175238 216732 175244
rect 216586 146024 216642 146033
rect 216586 145959 216642 145968
rect 216496 145716 216548 145722
rect 216496 145658 216548 145664
rect 216404 58608 216456 58614
rect 216404 58550 216456 58556
rect 216312 56432 216364 56438
rect 216312 56374 216364 56380
rect 216128 56024 216180 56030
rect 216128 55966 216180 55972
rect 216036 55956 216088 55962
rect 216036 55898 216088 55904
rect 215944 55140 215996 55146
rect 215944 55082 215996 55088
rect 214930 55040 214986 55049
rect 214930 54975 214986 54984
rect 214840 54596 214892 54602
rect 214840 54538 214892 54544
rect 216508 54534 216536 145658
rect 216600 59430 216628 145959
rect 216784 90001 216812 196959
rect 216876 145858 216904 270370
rect 216968 195265 216996 302087
rect 217048 268660 217100 268666
rect 217048 268602 217100 268608
rect 217060 268462 217088 268602
rect 217048 268456 217100 268462
rect 217048 268398 217100 268404
rect 216954 195256 217010 195265
rect 216954 195191 217010 195200
rect 216956 175228 217008 175234
rect 216956 175170 217008 175176
rect 216968 175137 216996 175170
rect 216954 175128 217010 175137
rect 216954 175063 217010 175072
rect 217060 162858 217088 268398
rect 217152 203017 217180 309975
rect 217244 270026 217272 375634
rect 217336 305017 217364 380734
rect 217520 377942 217548 480226
rect 217692 475380 217744 475386
rect 217692 475322 217744 475328
rect 217600 469124 217652 469130
rect 217600 469066 217652 469072
rect 217508 377936 217560 377942
rect 217414 377904 217470 377913
rect 217508 377878 217560 377884
rect 217414 377839 217470 377848
rect 217322 305008 217378 305017
rect 217322 304943 217378 304952
rect 217232 270020 217284 270026
rect 217232 269962 217284 269968
rect 217232 269068 217284 269074
rect 217232 269010 217284 269016
rect 217244 268705 217272 269010
rect 217230 268696 217286 268705
rect 217428 268666 217456 377839
rect 217612 376514 217640 469066
rect 217704 412049 217732 475322
rect 218060 467288 218112 467294
rect 218060 467230 218112 467236
rect 218072 466546 218100 467230
rect 218060 466540 218112 466546
rect 218060 466482 218112 466488
rect 217784 464568 217836 464574
rect 217784 464510 217836 464516
rect 217690 412040 217746 412049
rect 217690 411975 217746 411984
rect 217704 411369 217732 411975
rect 217690 411360 217746 411369
rect 217796 411330 217824 464510
rect 217968 422952 218020 422958
rect 217968 422894 218020 422900
rect 217980 416945 218008 422894
rect 217966 416936 218022 416945
rect 217966 416871 218022 416880
rect 217690 411295 217746 411304
rect 217784 411324 217836 411330
rect 217784 411266 217836 411272
rect 217874 409184 217930 409193
rect 217874 409119 217930 409128
rect 217888 379681 217916 409119
rect 217874 379672 217930 379681
rect 217784 379636 217836 379642
rect 217874 379607 217930 379616
rect 217784 379578 217836 379584
rect 217690 379536 217746 379545
rect 217690 379471 217746 379480
rect 217600 376508 217652 376514
rect 217600 376450 217652 376456
rect 217600 375828 217652 375834
rect 217600 375770 217652 375776
rect 217508 375352 217560 375358
rect 217508 375294 217560 375300
rect 217520 374921 217548 375294
rect 217506 374912 217562 374921
rect 217506 374847 217562 374856
rect 217612 354674 217640 375770
rect 217520 354646 217640 354674
rect 217520 311001 217548 354646
rect 217506 310992 217562 311001
rect 217562 310950 217640 310978
rect 217506 310927 217562 310936
rect 217506 307728 217562 307737
rect 217506 307663 217562 307672
rect 217520 306785 217548 307663
rect 217506 306776 217562 306785
rect 217506 306711 217562 306720
rect 217230 268631 217286 268640
rect 217416 268660 217468 268666
rect 217416 268602 217468 268608
rect 217414 203960 217470 203969
rect 217414 203895 217470 203904
rect 217138 203008 217194 203017
rect 217138 202943 217194 202952
rect 217230 198792 217286 198801
rect 217230 198727 217286 198736
rect 217048 162852 217100 162858
rect 217048 162794 217100 162800
rect 217048 145920 217100 145926
rect 217048 145862 217100 145868
rect 216864 145852 216916 145858
rect 216864 145794 216916 145800
rect 216956 145580 217008 145586
rect 216956 145522 217008 145528
rect 216968 144906 216996 145522
rect 216956 144900 217008 144906
rect 216956 144842 217008 144848
rect 216770 89992 216826 90001
rect 216770 89927 216826 89936
rect 216680 70372 216732 70378
rect 216680 70314 216732 70320
rect 216692 70009 216720 70314
rect 216678 70000 216734 70009
rect 216678 69935 216734 69944
rect 216678 68368 216734 68377
rect 216678 68303 216734 68312
rect 216692 67658 216720 68303
rect 216680 67652 216732 67658
rect 216680 67594 216732 67600
rect 216588 59424 216640 59430
rect 216588 59366 216640 59372
rect 217060 56098 217088 145862
rect 217140 144900 217192 144906
rect 217140 144842 217192 144848
rect 217048 56092 217100 56098
rect 217048 56034 217100 56040
rect 217152 54670 217180 144842
rect 217244 92857 217272 198727
rect 217324 162648 217376 162654
rect 217322 162616 217324 162625
rect 217376 162616 217378 162625
rect 217322 162551 217378 162560
rect 217428 96937 217456 203895
rect 217520 199889 217548 306711
rect 217612 203969 217640 310950
rect 217704 307873 217732 379471
rect 217690 307864 217746 307873
rect 217690 307799 217746 307808
rect 217598 203960 217654 203969
rect 217598 203895 217654 203904
rect 217598 203008 217654 203017
rect 217598 202943 217654 202952
rect 217506 199880 217562 199889
rect 217506 199815 217562 199824
rect 217520 198801 217548 199815
rect 217506 198792 217562 198801
rect 217506 198727 217562 198736
rect 217506 198112 217562 198121
rect 217506 198047 217562 198056
rect 217414 96928 217470 96937
rect 217414 96863 217470 96872
rect 217230 92848 217286 92857
rect 217230 92783 217286 92792
rect 217520 91089 217548 198047
rect 217612 95985 217640 202943
rect 217704 200841 217732 307799
rect 217796 303929 217824 379578
rect 217876 358284 217928 358290
rect 217876 358226 217928 358232
rect 217782 303920 217838 303929
rect 217782 303855 217838 303864
rect 217690 200832 217746 200841
rect 217690 200767 217746 200776
rect 217598 95976 217654 95985
rect 217598 95911 217654 95920
rect 217704 93809 217732 200767
rect 217796 197033 217824 303855
rect 217888 270366 217916 358226
rect 217980 310049 218008 416871
rect 218060 380044 218112 380050
rect 218060 379986 218112 379992
rect 218072 379642 218100 379986
rect 218060 379636 218112 379642
rect 218060 379578 218112 379584
rect 218164 375018 218192 485318
rect 218244 466540 218296 466546
rect 218244 466482 218296 466488
rect 218256 381546 218284 466482
rect 218244 381540 218296 381546
rect 218244 381482 218296 381488
rect 218348 379137 218376 488022
rect 219084 485178 219112 488022
rect 219176 485246 219204 488036
rect 219574 488022 219848 488050
rect 219164 485240 219216 485246
rect 219164 485182 219216 485188
rect 219072 485172 219124 485178
rect 219072 485114 219124 485120
rect 219716 485172 219768 485178
rect 219716 485114 219768 485120
rect 219164 484968 219216 484974
rect 219164 484910 219216 484916
rect 218704 478168 218756 478174
rect 218704 478110 218756 478116
rect 218334 379128 218390 379137
rect 218334 379063 218390 379072
rect 218348 378593 218376 379063
rect 218334 378584 218390 378593
rect 218334 378519 218390 378528
rect 218152 375012 218204 375018
rect 218152 374954 218204 374960
rect 218612 375012 218664 375018
rect 218612 374954 218664 374960
rect 218520 358760 218572 358766
rect 218520 358702 218572 358708
rect 217966 310040 218022 310049
rect 217966 309975 218022 309984
rect 217876 270360 217928 270366
rect 217876 270302 217928 270308
rect 217888 267734 217916 270302
rect 218428 270156 218480 270162
rect 218428 270098 218480 270104
rect 218152 269340 218204 269346
rect 218152 269282 218204 269288
rect 217888 267706 218008 267734
rect 217782 197024 217838 197033
rect 217782 196959 217838 196968
rect 217782 195256 217838 195265
rect 217782 195191 217838 195200
rect 217690 93800 217746 93809
rect 217690 93735 217746 93744
rect 217506 91080 217562 91089
rect 217506 91015 217562 91024
rect 217796 88233 217824 195191
rect 217876 162852 217928 162858
rect 217876 162794 217928 162800
rect 217888 161498 217916 162794
rect 217876 161492 217928 161498
rect 217876 161434 217928 161440
rect 217782 88224 217838 88233
rect 217782 88159 217838 88168
rect 217888 59566 217916 161434
rect 217980 146062 218008 267706
rect 217968 146056 218020 146062
rect 217968 145998 218020 146004
rect 218164 145790 218192 269282
rect 218440 268870 218468 270098
rect 218532 269550 218560 358702
rect 218624 270162 218652 374954
rect 218612 270156 218664 270162
rect 218612 270098 218664 270104
rect 218612 270020 218664 270026
rect 218612 269962 218664 269968
rect 218520 269544 218572 269550
rect 218520 269486 218572 269492
rect 218624 269414 218652 269962
rect 218612 269408 218664 269414
rect 218612 269350 218664 269356
rect 218428 268864 218480 268870
rect 218428 268806 218480 268812
rect 218520 268796 218572 268802
rect 218520 268738 218572 268744
rect 218532 268530 218560 268738
rect 218520 268524 218572 268530
rect 218520 268466 218572 268472
rect 218242 165608 218298 165617
rect 218242 165543 218298 165552
rect 218152 145784 218204 145790
rect 218152 145726 218204 145732
rect 217966 68368 218022 68377
rect 217966 68303 218022 68312
rect 217876 59560 217928 59566
rect 217876 59502 217928 59508
rect 217980 59362 218008 68303
rect 217968 59356 218020 59362
rect 217968 59298 218020 59304
rect 218256 57798 218284 165543
rect 218336 164144 218388 164150
rect 218336 164086 218388 164092
rect 218244 57792 218296 57798
rect 218244 57734 218296 57740
rect 218348 54942 218376 164086
rect 218532 162858 218560 268466
rect 218612 252544 218664 252550
rect 218612 252486 218664 252492
rect 218520 162852 218572 162858
rect 218520 162794 218572 162800
rect 218624 146169 218652 252486
rect 218610 146160 218666 146169
rect 218610 146095 218666 146104
rect 218428 145988 218480 145994
rect 218428 145930 218480 145936
rect 218336 54936 218388 54942
rect 218336 54878 218388 54884
rect 218440 54806 218468 145930
rect 218520 145512 218572 145518
rect 218520 145454 218572 145460
rect 218532 59702 218560 145454
rect 218520 59696 218572 59702
rect 218520 59638 218572 59644
rect 218624 56234 218652 146095
rect 218716 57254 218744 478110
rect 219072 475584 219124 475590
rect 219072 475526 219124 475532
rect 218796 474156 218848 474162
rect 218796 474098 218848 474104
rect 218808 57390 218836 474098
rect 218888 467220 218940 467226
rect 218888 467162 218940 467168
rect 218900 165102 218928 467162
rect 218978 465760 219034 465769
rect 218978 465695 219034 465704
rect 218992 165238 219020 465695
rect 219084 271454 219112 475526
rect 219176 378826 219204 484910
rect 219532 484220 219584 484226
rect 219532 484162 219584 484168
rect 219256 411324 219308 411330
rect 219256 411266 219308 411272
rect 219164 378820 219216 378826
rect 219164 378762 219216 378768
rect 219268 376242 219296 411266
rect 219544 382430 219572 484162
rect 219624 484152 219676 484158
rect 219624 484094 219676 484100
rect 219636 417450 219664 484094
rect 219624 417444 219676 417450
rect 219624 417386 219676 417392
rect 219532 382424 219584 382430
rect 219532 382366 219584 382372
rect 219532 382288 219584 382294
rect 219532 382230 219584 382236
rect 219440 379704 219492 379710
rect 219440 379646 219492 379652
rect 219348 377528 219400 377534
rect 219348 377470 219400 377476
rect 219256 376236 219308 376242
rect 219256 376178 219308 376184
rect 219256 374672 219308 374678
rect 219256 374614 219308 374620
rect 219164 358556 219216 358562
rect 219164 358498 219216 358504
rect 219072 271448 219124 271454
rect 219072 271390 219124 271396
rect 219070 269920 219126 269929
rect 219070 269855 219072 269864
rect 219124 269855 219126 269864
rect 219072 269826 219124 269832
rect 219084 269498 219112 269826
rect 219176 269618 219204 358498
rect 219268 273562 219296 374614
rect 219256 273556 219308 273562
rect 219256 273498 219308 273504
rect 219360 269958 219388 377470
rect 219348 269952 219400 269958
rect 219348 269894 219400 269900
rect 219164 269612 219216 269618
rect 219164 269554 219216 269560
rect 219256 269544 219308 269550
rect 219084 269470 219204 269498
rect 219256 269486 219308 269492
rect 219072 269408 219124 269414
rect 219072 269350 219124 269356
rect 218980 165232 219032 165238
rect 218980 165174 219032 165180
rect 218888 165096 218940 165102
rect 218888 165038 218940 165044
rect 219084 164150 219112 269350
rect 219072 164144 219124 164150
rect 219072 164086 219124 164092
rect 218980 162852 219032 162858
rect 218980 162794 219032 162800
rect 218992 161566 219020 162794
rect 219176 161838 219204 269470
rect 219164 161832 219216 161838
rect 219164 161774 219216 161780
rect 218980 161560 219032 161566
rect 218980 161502 219032 161508
rect 218888 145784 218940 145790
rect 218888 145726 218940 145732
rect 218796 57384 218848 57390
rect 218796 57326 218848 57332
rect 218704 57248 218756 57254
rect 218704 57190 218756 57196
rect 218612 56228 218664 56234
rect 218612 56170 218664 56176
rect 218900 55214 218928 145726
rect 218992 59498 219020 161502
rect 219268 146130 219296 269486
rect 219360 269142 219388 269894
rect 219348 269136 219400 269142
rect 219348 269078 219400 269084
rect 219452 269006 219480 379646
rect 219544 376038 219572 382230
rect 219728 379370 219756 485114
rect 219820 379506 219848 488022
rect 219912 488022 220018 488050
rect 220096 488022 220478 488050
rect 219912 484226 219940 488022
rect 219992 484424 220044 484430
rect 219992 484366 220044 484372
rect 219900 484220 219952 484226
rect 219900 484162 219952 484168
rect 219900 382424 219952 382430
rect 219900 382366 219952 382372
rect 219808 379500 219860 379506
rect 219808 379442 219860 379448
rect 219624 379364 219676 379370
rect 219624 379306 219676 379312
rect 219716 379364 219768 379370
rect 219716 379306 219768 379312
rect 219636 378554 219664 379306
rect 219808 379228 219860 379234
rect 219808 379170 219860 379176
rect 219716 378956 219768 378962
rect 219716 378898 219768 378904
rect 219728 378758 219756 378898
rect 219716 378752 219768 378758
rect 219716 378694 219768 378700
rect 219624 378548 219676 378554
rect 219624 378490 219676 378496
rect 219532 376032 219584 376038
rect 219532 375974 219584 375980
rect 219636 269278 219664 378490
rect 219820 270502 219848 379170
rect 219912 379166 219940 382366
rect 219900 379160 219952 379166
rect 219900 379102 219952 379108
rect 219900 378752 219952 378758
rect 219900 378694 219952 378700
rect 219808 270496 219860 270502
rect 219808 270438 219860 270444
rect 219912 270434 219940 378694
rect 219900 270428 219952 270434
rect 219900 270370 219952 270376
rect 219716 270088 219768 270094
rect 219716 270030 219768 270036
rect 219624 269272 219676 269278
rect 219624 269214 219676 269220
rect 219624 269136 219676 269142
rect 219624 269078 219676 269084
rect 219440 269000 219492 269006
rect 219440 268942 219492 268948
rect 219452 262954 219480 268942
rect 219440 262948 219492 262954
rect 219440 262890 219492 262896
rect 219636 164218 219664 269078
rect 219728 267734 219756 270030
rect 219900 269612 219952 269618
rect 219900 269554 219952 269560
rect 219728 267706 219848 267734
rect 219716 262948 219768 262954
rect 219716 262890 219768 262896
rect 219624 164212 219676 164218
rect 219624 164154 219676 164160
rect 219348 162784 219400 162790
rect 219348 162726 219400 162732
rect 219360 162450 219388 162726
rect 219348 162444 219400 162450
rect 219348 162386 219400 162392
rect 219532 161832 219584 161838
rect 219532 161774 219584 161780
rect 219256 146124 219308 146130
rect 219256 146066 219308 146072
rect 219070 60616 219126 60625
rect 219070 60551 219126 60560
rect 218980 59492 219032 59498
rect 218980 59434 219032 59440
rect 219084 58682 219112 60551
rect 219072 58676 219124 58682
rect 219072 58618 219124 58624
rect 218888 55208 218940 55214
rect 218888 55150 218940 55156
rect 218428 54800 218480 54806
rect 218428 54742 218480 54748
rect 219268 54738 219296 146066
rect 219544 55078 219572 161774
rect 219532 55072 219584 55078
rect 219532 55014 219584 55020
rect 219636 55010 219664 164154
rect 219728 145450 219756 262890
rect 219820 145994 219848 267706
rect 219912 145994 219940 269554
rect 219808 145988 219860 145994
rect 219808 145930 219860 145936
rect 219900 145988 219952 145994
rect 219900 145930 219952 145936
rect 219716 145444 219768 145450
rect 219716 145386 219768 145392
rect 219624 55004 219676 55010
rect 219624 54946 219676 54952
rect 219728 54874 219756 145386
rect 219820 145382 219848 145930
rect 219898 145888 219954 145897
rect 219898 145823 219954 145832
rect 219808 145376 219860 145382
rect 219808 145318 219860 145324
rect 219912 56302 219940 145823
rect 220004 56574 220032 484366
rect 220096 484158 220124 488022
rect 220084 484152 220136 484158
rect 220084 484094 220136 484100
rect 220924 465730 220952 488036
rect 221016 488022 221398 488050
rect 221016 466410 221044 488022
rect 221752 485110 221780 488036
rect 222242 488022 222608 488050
rect 221740 485104 221792 485110
rect 221740 485046 221792 485052
rect 222580 482361 222608 488022
rect 222672 484430 222700 488036
rect 223162 488022 223528 488050
rect 223622 488022 223712 488050
rect 223990 488022 224080 488050
rect 223500 485110 223528 488022
rect 223488 485104 223540 485110
rect 223488 485046 223540 485052
rect 222660 484424 222712 484430
rect 222660 484366 222712 484372
rect 223580 483404 223632 483410
rect 223580 483346 223632 483352
rect 222566 482352 222622 482361
rect 222566 482287 222622 482296
rect 223592 474065 223620 483346
rect 223684 478281 223712 488022
rect 224052 485178 224080 488022
rect 224144 488022 224434 488050
rect 224040 485172 224092 485178
rect 224040 485114 224092 485120
rect 224144 483410 224172 488022
rect 224880 484537 224908 488036
rect 225370 488022 225644 488050
rect 225616 485246 225644 488022
rect 225604 485240 225656 485246
rect 225708 485217 225736 488036
rect 225604 485182 225656 485188
rect 225694 485208 225750 485217
rect 225694 485143 225750 485152
rect 226168 485081 226196 488036
rect 226154 485072 226210 485081
rect 226154 485007 226210 485016
rect 224866 484528 224922 484537
rect 224866 484463 224922 484472
rect 226628 484294 226656 488036
rect 226720 488022 227102 488050
rect 227272 488022 227562 488050
rect 226616 484288 226668 484294
rect 226616 484230 226668 484236
rect 226720 484140 226748 488022
rect 226352 484112 226748 484140
rect 224132 483404 224184 483410
rect 224132 483346 224184 483352
rect 223670 478272 223726 478281
rect 223670 478207 223726 478216
rect 223578 474056 223634 474065
rect 223578 473991 223634 474000
rect 226352 472802 226380 484112
rect 226340 472796 226392 472802
rect 226340 472738 226392 472744
rect 227272 472666 227300 488022
rect 227628 484288 227680 484294
rect 227628 484230 227680 484236
rect 227640 483682 227668 484230
rect 227720 484152 227772 484158
rect 227720 484094 227772 484100
rect 227628 483676 227680 483682
rect 227628 483618 227680 483624
rect 227732 474473 227760 484094
rect 227916 483750 227944 488036
rect 228008 488022 228390 488050
rect 228560 488022 228850 488050
rect 229204 488022 229310 488050
rect 229480 488022 229770 488050
rect 230154 488022 230428 488050
rect 230614 488022 230704 488050
rect 227904 483744 227956 483750
rect 227904 483686 227956 483692
rect 228008 476921 228036 488022
rect 228560 484158 228588 488022
rect 228548 484152 228600 484158
rect 228548 484094 228600 484100
rect 229100 484152 229152 484158
rect 229100 484094 229152 484100
rect 227994 476912 228050 476921
rect 227994 476847 228050 476856
rect 227718 474464 227774 474473
rect 227718 474399 227774 474408
rect 227260 472660 227312 472666
rect 227260 472602 227312 472608
rect 229112 472569 229140 484094
rect 229204 475386 229232 488022
rect 229480 484158 229508 488022
rect 229468 484152 229520 484158
rect 229468 484094 229520 484100
rect 230400 483721 230428 488022
rect 230676 485625 230704 488022
rect 230768 488022 231058 488050
rect 231534 488022 231808 488050
rect 231902 488022 232176 488050
rect 230662 485616 230718 485625
rect 230662 485551 230718 485560
rect 230386 483712 230442 483721
rect 230386 483647 230442 483656
rect 229192 475380 229244 475386
rect 229192 475322 229244 475328
rect 230768 474201 230796 488022
rect 231780 485081 231808 488022
rect 231766 485072 231822 485081
rect 231766 485007 231822 485016
rect 232148 480865 232176 488022
rect 232332 485217 232360 488036
rect 232424 488022 232806 488050
rect 232318 485208 232374 485217
rect 232318 485143 232374 485152
rect 232134 480856 232190 480865
rect 232134 480791 232190 480800
rect 232424 475522 232452 488022
rect 233252 485314 233280 488036
rect 233344 488022 233726 488050
rect 234110 488022 234384 488050
rect 233240 485308 233292 485314
rect 233240 485250 233292 485256
rect 233344 479641 233372 488022
rect 234356 485489 234384 488022
rect 234342 485480 234398 485489
rect 234342 485415 234398 485424
rect 234540 485382 234568 488036
rect 234632 488022 235014 488050
rect 235490 488022 235856 488050
rect 234528 485376 234580 485382
rect 234528 485318 234580 485324
rect 233330 479632 233386 479641
rect 233330 479567 233386 479576
rect 234632 476785 234660 488022
rect 235828 485761 235856 488022
rect 235814 485752 235870 485761
rect 235814 485687 235870 485696
rect 235920 485353 235948 488036
rect 236318 488022 236408 488050
rect 235906 485344 235962 485353
rect 235906 485279 235962 485288
rect 236000 484152 236052 484158
rect 236000 484094 236052 484100
rect 234618 476776 234674 476785
rect 234618 476711 234674 476720
rect 232412 475516 232464 475522
rect 232412 475458 232464 475464
rect 230754 474192 230810 474201
rect 230754 474127 230810 474136
rect 229098 472560 229154 472569
rect 229098 472495 229154 472504
rect 221004 466404 221056 466410
rect 221004 466346 221056 466352
rect 236012 465798 236040 484094
rect 236380 482497 236408 488022
rect 236472 488022 236762 488050
rect 236840 488022 237222 488050
rect 237392 488022 237682 488050
rect 237760 488022 238142 488050
rect 238220 488022 238510 488050
rect 238772 488022 238970 488050
rect 239446 488022 239720 488050
rect 239906 488022 240088 488050
rect 236366 482488 236422 482497
rect 236366 482423 236422 482432
rect 236472 475590 236500 488022
rect 236840 484158 236868 488022
rect 236828 484152 236880 484158
rect 236828 484094 236880 484100
rect 236460 475584 236512 475590
rect 236460 475526 236512 475532
rect 237392 472734 237420 488022
rect 237760 484106 237788 488022
rect 237484 484078 237788 484106
rect 237484 475454 237512 484078
rect 238220 478310 238248 488022
rect 238208 478304 238260 478310
rect 238208 478246 238260 478252
rect 238772 478174 238800 488022
rect 239692 485450 239720 488022
rect 240060 485518 240088 488022
rect 240152 488022 240258 488050
rect 240336 488022 240718 488050
rect 240796 488022 241178 488050
rect 240048 485512 240100 485518
rect 240048 485454 240100 485460
rect 239680 485444 239732 485450
rect 239680 485386 239732 485392
rect 238760 478168 238812 478174
rect 238760 478110 238812 478116
rect 237472 475448 237524 475454
rect 237472 475390 237524 475396
rect 240152 474094 240180 488022
rect 240336 484140 240364 488022
rect 240244 484112 240364 484140
rect 240244 474337 240272 484112
rect 240230 474328 240286 474337
rect 240230 474263 240286 474272
rect 240140 474088 240192 474094
rect 240140 474030 240192 474036
rect 240796 474026 240824 488022
rect 241520 484152 241572 484158
rect 241520 484094 241572 484100
rect 240784 474020 240836 474026
rect 240784 473962 240836 473968
rect 237380 472728 237432 472734
rect 237380 472670 237432 472676
rect 241532 465934 241560 484094
rect 241624 472870 241652 488036
rect 242084 485586 242112 488036
rect 242176 488022 242466 488050
rect 242942 488022 243032 488050
rect 242072 485580 242124 485586
rect 242072 485522 242124 485528
rect 242176 484158 242204 488022
rect 242164 484152 242216 484158
rect 242164 484094 242216 484100
rect 242900 482588 242952 482594
rect 242900 482530 242952 482536
rect 241612 472864 241664 472870
rect 241612 472806 241664 472812
rect 241520 465928 241572 465934
rect 241520 465870 241572 465876
rect 236000 465792 236052 465798
rect 236000 465734 236052 465740
rect 242912 465730 242940 482530
rect 243004 479602 243032 488022
rect 243096 488022 243386 488050
rect 243862 488022 244136 488050
rect 244322 488022 244504 488050
rect 243096 482594 243124 488022
rect 243084 482588 243136 482594
rect 243084 482530 243136 482536
rect 244108 481098 244136 488022
rect 244096 481092 244148 481098
rect 244096 481034 244148 481040
rect 242992 479596 243044 479602
rect 242992 479538 243044 479544
rect 244476 476814 244504 488022
rect 244660 482390 244688 488036
rect 244752 488022 245134 488050
rect 245304 488022 245594 488050
rect 244648 482384 244700 482390
rect 244648 482326 244700 482332
rect 244464 476808 244516 476814
rect 244464 476750 244516 476756
rect 244752 476626 244780 488022
rect 244292 476598 244780 476626
rect 244292 465866 244320 476598
rect 245304 476114 245332 488022
rect 246040 483818 246068 488036
rect 246132 488022 246422 488050
rect 246500 488022 246882 488050
rect 246028 483812 246080 483818
rect 246028 483754 246080 483760
rect 246132 476882 246160 488022
rect 246500 479534 246528 488022
rect 247328 481001 247356 488036
rect 247420 488022 247802 488050
rect 248278 488022 248368 488050
rect 248646 488022 248736 488050
rect 247314 480992 247370 481001
rect 247314 480927 247370 480936
rect 246488 479528 246540 479534
rect 246488 479470 246540 479476
rect 247420 478378 247448 488022
rect 248340 482322 248368 488022
rect 248708 484945 248736 488022
rect 248800 488022 249090 488050
rect 249168 488022 249550 488050
rect 248694 484936 248750 484945
rect 248694 484871 248750 484880
rect 248328 482316 248380 482322
rect 248328 482258 248380 482264
rect 248420 480888 248472 480894
rect 248420 480830 248472 480836
rect 247408 478372 247460 478378
rect 247408 478314 247460 478320
rect 246120 476876 246172 476882
rect 246120 476818 246172 476824
rect 244384 476086 245332 476114
rect 244384 474162 244412 476086
rect 244372 474156 244424 474162
rect 244372 474098 244424 474104
rect 248432 466070 248460 480830
rect 248800 470594 248828 488022
rect 249168 480894 249196 488022
rect 249156 480888 249208 480894
rect 249156 480830 249208 480836
rect 249892 480888 249944 480894
rect 249892 480830 249944 480836
rect 249800 478236 249852 478242
rect 249800 478178 249852 478184
rect 248524 470566 248828 470594
rect 248524 466138 248552 470566
rect 249812 466206 249840 478178
rect 249904 468518 249932 480830
rect 249996 468586 250024 488036
rect 250088 488022 250470 488050
rect 250548 488022 250838 488050
rect 251314 488022 251404 488050
rect 250088 480894 250116 488022
rect 250076 480888 250128 480894
rect 250076 480830 250128 480836
rect 250548 478242 250576 488022
rect 251376 481166 251404 488022
rect 251468 488022 251758 488050
rect 251928 488022 252218 488050
rect 252602 488022 252968 488050
rect 253062 488022 253152 488050
rect 251364 481160 251416 481166
rect 251364 481102 251416 481108
rect 251180 480888 251232 480894
rect 251180 480830 251232 480836
rect 250536 478236 250588 478242
rect 250536 478178 250588 478184
rect 249984 468580 250036 468586
rect 249984 468522 250036 468528
rect 249892 468512 249944 468518
rect 249892 468454 249944 468460
rect 251192 467158 251220 480830
rect 251468 478122 251496 488022
rect 251548 481160 251600 481166
rect 251548 481102 251600 481108
rect 251284 478094 251496 478122
rect 251284 467362 251312 478094
rect 251560 473354 251588 481102
rect 251928 480894 251956 488022
rect 252940 483857 252968 488022
rect 252926 483848 252982 483857
rect 252926 483783 252982 483792
rect 253124 481030 253152 488022
rect 253216 488022 253506 488050
rect 253982 488022 254072 488050
rect 253112 481024 253164 481030
rect 253112 480966 253164 480972
rect 251916 480888 251968 480894
rect 251916 480830 251968 480836
rect 253216 479670 253244 488022
rect 253940 480888 253992 480894
rect 253940 480830 253992 480836
rect 253204 479664 253256 479670
rect 253204 479606 253256 479612
rect 251376 473326 251588 473354
rect 251376 471306 251404 473326
rect 251364 471300 251416 471306
rect 251364 471242 251416 471248
rect 251272 467356 251324 467362
rect 251272 467298 251324 467304
rect 251180 467152 251232 467158
rect 251180 467094 251232 467100
rect 249800 466200 249852 466206
rect 249800 466142 249852 466148
rect 248512 466132 248564 466138
rect 248512 466074 248564 466080
rect 248420 466064 248472 466070
rect 248420 466006 248472 466012
rect 253952 466002 253980 480830
rect 254044 468722 254072 488022
rect 254136 488022 254426 488050
rect 254504 488022 254794 488050
rect 254136 480894 254164 488022
rect 254124 480888 254176 480894
rect 254124 480830 254176 480836
rect 254504 479738 254532 488022
rect 255240 482458 255268 488036
rect 255332 488022 255714 488050
rect 255792 488022 256174 488050
rect 256344 488022 256634 488050
rect 256712 488022 257002 488050
rect 257478 488022 257568 488050
rect 255228 482452 255280 482458
rect 255228 482394 255280 482400
rect 254492 479732 254544 479738
rect 254492 479674 254544 479680
rect 255332 468790 255360 488022
rect 255792 476114 255820 488022
rect 255424 476086 255820 476114
rect 255424 471374 255452 476086
rect 256344 475425 256372 488022
rect 256330 475416 256386 475425
rect 256330 475351 256386 475360
rect 255412 471368 255464 471374
rect 255412 471310 255464 471316
rect 255320 468784 255372 468790
rect 255320 468726 255372 468732
rect 254032 468716 254084 468722
rect 254032 468658 254084 468664
rect 256712 467430 256740 488022
rect 257540 482594 257568 488022
rect 257632 488022 257922 488050
rect 258092 488022 258382 488050
rect 258552 488022 258842 488050
rect 258920 488022 259210 488050
rect 259472 488022 259670 488050
rect 259748 488022 260130 488050
rect 260208 488022 260590 488050
rect 257528 482588 257580 482594
rect 257528 482530 257580 482536
rect 257632 474298 257660 488022
rect 257620 474292 257672 474298
rect 257620 474234 257672 474240
rect 256700 467424 256752 467430
rect 256700 467366 256752 467372
rect 258092 467226 258120 488022
rect 258552 476950 258580 488022
rect 258540 476944 258592 476950
rect 258540 476886 258592 476892
rect 258920 476114 258948 488022
rect 258184 476086 258948 476114
rect 258184 472938 258212 476086
rect 259472 475658 259500 488022
rect 259748 477018 259776 488022
rect 260208 478378 260236 488022
rect 260944 479874 260972 488036
rect 261404 482526 261432 488036
rect 261496 488022 261878 488050
rect 262232 488022 262338 488050
rect 262508 488022 262798 488050
rect 262876 488022 263166 488050
rect 261392 482520 261444 482526
rect 261392 482462 261444 482468
rect 260932 479868 260984 479874
rect 260932 479810 260984 479816
rect 260196 478372 260248 478378
rect 260196 478314 260248 478320
rect 259736 477012 259788 477018
rect 259736 476954 259788 476960
rect 261496 476114 261524 488022
rect 262232 481234 262260 488022
rect 262508 485774 262536 488022
rect 262324 485746 262536 485774
rect 262220 481228 262272 481234
rect 262220 481170 262272 481176
rect 262324 480978 262352 485746
rect 262588 481228 262640 481234
rect 262588 481170 262640 481176
rect 260852 476086 261524 476114
rect 262232 480950 262352 480978
rect 259460 475652 259512 475658
rect 259460 475594 259512 475600
rect 258172 472932 258224 472938
rect 258172 472874 258224 472880
rect 260852 467294 260880 476086
rect 260840 467288 260892 467294
rect 260840 467230 260892 467236
rect 258080 467220 258132 467226
rect 258080 467162 258132 467168
rect 262232 466274 262260 480950
rect 262312 480888 262364 480894
rect 262312 480830 262364 480836
rect 262324 473006 262352 480830
rect 262600 476114 262628 481170
rect 262876 480894 262904 488022
rect 262864 480888 262916 480894
rect 262864 480830 262916 480836
rect 263612 477154 263640 488036
rect 263704 488022 264086 488050
rect 264256 488022 264546 488050
rect 265022 488022 265296 488050
rect 263600 477148 263652 477154
rect 263600 477090 263652 477096
rect 263704 477086 263732 488022
rect 264256 477222 264284 488022
rect 265164 484220 265216 484226
rect 265164 484162 265216 484168
rect 265072 484152 265124 484158
rect 265072 484094 265124 484100
rect 264980 484084 265032 484090
rect 264980 484026 265032 484032
rect 264244 477216 264296 477222
rect 264244 477158 264296 477164
rect 263692 477080 263744 477086
rect 263692 477022 263744 477028
rect 262416 476086 262628 476114
rect 262416 474230 262444 476086
rect 262404 474224 262456 474230
rect 262404 474166 262456 474172
rect 262312 473000 262364 473006
rect 262312 472942 262364 472948
rect 264992 466410 265020 484026
rect 265084 468489 265112 484094
rect 265176 468994 265204 484162
rect 265268 479806 265296 488022
rect 265360 484090 265388 488036
rect 265544 488022 265834 488050
rect 265912 488022 266294 488050
rect 266556 488022 266754 488050
rect 266832 488022 267122 488050
rect 267200 488022 267582 488050
rect 265544 484158 265572 488022
rect 265912 484226 265940 488022
rect 265900 484220 265952 484226
rect 265900 484162 265952 484168
rect 266452 484220 266504 484226
rect 266452 484162 266504 484168
rect 265532 484152 265584 484158
rect 265532 484094 265584 484100
rect 266360 484152 266412 484158
rect 266360 484094 266412 484100
rect 265348 484084 265400 484090
rect 265348 484026 265400 484032
rect 265256 479800 265308 479806
rect 265256 479742 265308 479748
rect 266372 469198 266400 484094
rect 266360 469192 266412 469198
rect 266360 469134 266412 469140
rect 265164 468988 265216 468994
rect 265164 468930 265216 468936
rect 266464 468654 266492 484162
rect 266556 469062 266584 488022
rect 266832 484158 266860 488022
rect 267200 484226 267228 488022
rect 267188 484220 267240 484226
rect 267188 484162 267240 484168
rect 266820 484152 266872 484158
rect 266820 484094 266872 484100
rect 268028 483886 268056 488036
rect 268120 488022 268502 488050
rect 268978 488022 269068 488050
rect 268016 483880 268068 483886
rect 268016 483822 268068 483828
rect 268120 470594 268148 488022
rect 269040 483954 269068 488022
rect 269132 488022 269330 488050
rect 269806 488022 270080 488050
rect 270266 488022 270448 488050
rect 269028 483948 269080 483954
rect 269028 483890 269080 483896
rect 267752 470566 268148 470594
rect 266544 469056 266596 469062
rect 266544 468998 266596 469004
rect 267752 468858 267780 470566
rect 267740 468852 267792 468858
rect 267740 468794 267792 468800
rect 266452 468648 266504 468654
rect 266452 468590 266504 468596
rect 265070 468480 265126 468489
rect 265070 468415 265126 468424
rect 264980 466404 265032 466410
rect 264980 466346 265032 466352
rect 269132 466342 269160 488022
rect 270052 481302 270080 488022
rect 270040 481296 270092 481302
rect 270040 481238 270092 481244
rect 270420 481234 270448 488022
rect 270512 488022 270710 488050
rect 270880 488022 271170 488050
rect 271554 488022 271828 488050
rect 270408 481228 270460 481234
rect 270408 481170 270460 481176
rect 270512 470082 270540 488022
rect 270880 475794 270908 488022
rect 271800 481166 271828 488022
rect 271892 488022 271998 488050
rect 271788 481160 271840 481166
rect 271788 481102 271840 481108
rect 270868 475788 270920 475794
rect 270868 475730 270920 475736
rect 270500 470076 270552 470082
rect 270500 470018 270552 470024
rect 269120 466336 269172 466342
rect 269120 466278 269172 466284
rect 262220 466268 262272 466274
rect 262220 466210 262272 466216
rect 253940 465996 253992 466002
rect 253940 465938 253992 465944
rect 244280 465860 244332 465866
rect 244280 465802 244332 465808
rect 220912 465724 220964 465730
rect 220912 465666 220964 465672
rect 242900 465724 242952 465730
rect 242900 465666 242952 465672
rect 271892 464370 271920 488022
rect 272444 482662 272472 488036
rect 272536 488022 272918 488050
rect 272432 482656 272484 482662
rect 272432 482598 272484 482604
rect 272536 470594 272564 488022
rect 271984 470566 272564 470594
rect 271984 469130 272012 470566
rect 271972 469124 272024 469130
rect 271972 469066 272024 469072
rect 273272 467498 273300 488036
rect 273456 488022 273746 488050
rect 273824 488022 274206 488050
rect 274682 488022 274772 488050
rect 273352 477896 273404 477902
rect 273352 477838 273404 477844
rect 273364 473074 273392 477838
rect 273456 474366 273484 488022
rect 273824 477902 273852 488022
rect 273812 477896 273864 477902
rect 273812 477838 273864 477844
rect 274744 477290 274772 488022
rect 274836 488022 275126 488050
rect 275204 488022 275494 488050
rect 275664 488022 275954 488050
rect 276032 488022 276414 488050
rect 276584 488022 276874 488050
rect 276952 488022 277334 488050
rect 277504 488022 277702 488050
rect 277872 488022 278162 488050
rect 278638 488022 278728 488050
rect 274732 477284 274784 477290
rect 274732 477226 274784 477232
rect 274836 476114 274864 488022
rect 275204 479942 275232 488022
rect 275192 479936 275244 479942
rect 275192 479878 275244 479884
rect 275664 478446 275692 488022
rect 275652 478440 275704 478446
rect 275652 478382 275704 478388
rect 274652 476086 274864 476114
rect 274652 475726 274680 476086
rect 274640 475720 274692 475726
rect 274640 475662 274692 475668
rect 273444 474360 273496 474366
rect 273444 474302 273496 474308
rect 273352 473068 273404 473074
rect 273352 473010 273404 473016
rect 276032 468926 276060 488022
rect 276584 477358 276612 488022
rect 276572 477352 276624 477358
rect 276572 477294 276624 477300
rect 276952 476114 276980 488022
rect 277400 477896 277452 477902
rect 277400 477838 277452 477844
rect 276124 476086 276980 476114
rect 276124 474609 276152 476086
rect 276110 474600 276166 474609
rect 276110 474535 276166 474544
rect 276020 468920 276072 468926
rect 276020 468862 276072 468868
rect 273260 467492 273312 467498
rect 273260 467434 273312 467440
rect 277412 465662 277440 477838
rect 277504 467566 277532 488022
rect 277872 477902 277900 488022
rect 278700 482730 278728 488022
rect 278884 488022 279082 488050
rect 279160 488022 279542 488050
rect 279926 488022 280108 488050
rect 278688 482724 278740 482730
rect 278688 482666 278740 482672
rect 278884 480010 278912 488022
rect 278872 480004 278924 480010
rect 278872 479946 278924 479952
rect 277860 477896 277912 477902
rect 277860 477838 277912 477844
rect 279160 476114 279188 488022
rect 280080 482798 280108 488022
rect 280172 488022 280370 488050
rect 280846 488022 281120 488050
rect 281306 488022 281488 488050
rect 281674 488022 281764 488050
rect 280068 482792 280120 482798
rect 280068 482734 280120 482740
rect 278792 476086 279188 476114
rect 278792 475862 278820 476086
rect 278780 475856 278832 475862
rect 278780 475798 278832 475804
rect 280172 473142 280200 488022
rect 281092 483993 281120 488022
rect 281460 484090 281488 488022
rect 281448 484084 281500 484090
rect 281448 484026 281500 484032
rect 281078 483984 281134 483993
rect 281078 483919 281134 483928
rect 281736 480146 281764 488022
rect 281828 488022 282118 488050
rect 282288 488022 282578 488050
rect 282932 488022 283038 488050
rect 283116 488022 283498 488050
rect 283576 488022 283866 488050
rect 284342 488022 284432 488050
rect 281724 480140 281776 480146
rect 281724 480082 281776 480088
rect 281828 480026 281856 488022
rect 281552 479998 281856 480026
rect 280160 473136 280212 473142
rect 280160 473078 280212 473084
rect 281552 470150 281580 479998
rect 282288 476114 282316 488022
rect 281644 476086 282316 476114
rect 281540 470144 281592 470150
rect 281540 470086 281592 470092
rect 281644 469878 281672 476086
rect 282932 470422 282960 488022
rect 283116 484140 283144 488022
rect 283024 484112 283144 484140
rect 282920 470416 282972 470422
rect 282920 470358 282972 470364
rect 283024 470354 283052 484112
rect 283576 470594 283604 488022
rect 284300 484152 284352 484158
rect 284300 484094 284352 484100
rect 283116 470566 283604 470594
rect 283116 470490 283144 470566
rect 283104 470484 283156 470490
rect 283104 470426 283156 470432
rect 283012 470348 283064 470354
rect 283012 470290 283064 470296
rect 284312 469946 284340 484094
rect 284404 470014 284432 488022
rect 284772 482866 284800 488036
rect 284864 488022 285246 488050
rect 284864 484158 284892 488022
rect 284852 484152 284904 484158
rect 284852 484094 284904 484100
rect 284760 482860 284812 482866
rect 284760 482802 284812 482808
rect 284392 470008 284444 470014
rect 284392 469950 284444 469956
rect 284300 469940 284352 469946
rect 284300 469882 284352 469888
rect 281632 469872 281684 469878
rect 281632 469814 281684 469820
rect 277492 467560 277544 467566
rect 277492 467502 277544 467508
rect 277400 465656 277452 465662
rect 277400 465598 277452 465604
rect 285692 465594 285720 488036
rect 285784 488022 286074 488050
rect 286152 488022 286534 488050
rect 285784 470218 285812 488022
rect 286152 471510 286180 488022
rect 286980 484090 287008 488036
rect 287164 488022 287454 488050
rect 287532 488022 287822 488050
rect 287992 488022 288282 488050
rect 288452 488022 288742 488050
rect 288912 488022 289202 488050
rect 289678 488022 289768 488050
rect 287060 484152 287112 484158
rect 287060 484094 287112 484100
rect 286968 484084 287020 484090
rect 286968 484026 287020 484032
rect 286140 471504 286192 471510
rect 286140 471446 286192 471452
rect 287072 470286 287100 484094
rect 287164 471442 287192 488022
rect 287152 471436 287204 471442
rect 287152 471378 287204 471384
rect 287532 471238 287560 488022
rect 287992 484158 288020 488022
rect 287980 484152 288032 484158
rect 287980 484094 288032 484100
rect 288452 471782 288480 488022
rect 288912 478582 288940 488022
rect 289740 481370 289768 488022
rect 289832 488022 290030 488050
rect 290200 488022 290490 488050
rect 290568 488022 290950 488050
rect 291212 488022 291410 488050
rect 291488 488022 291870 488050
rect 291948 488022 292238 488050
rect 292714 488022 292804 488050
rect 289728 481364 289780 481370
rect 289728 481306 289780 481312
rect 288900 478576 288952 478582
rect 288900 478518 288952 478524
rect 288440 471776 288492 471782
rect 288440 471718 288492 471724
rect 287520 471232 287572 471238
rect 287520 471174 287572 471180
rect 289832 470558 289860 488022
rect 289912 484152 289964 484158
rect 289912 484094 289964 484100
rect 289924 474502 289952 484094
rect 289912 474496 289964 474502
rect 289912 474438 289964 474444
rect 290200 474434 290228 488022
rect 290568 484158 290596 488022
rect 290556 484152 290608 484158
rect 290556 484094 290608 484100
rect 290188 474428 290240 474434
rect 290188 474370 290240 474376
rect 291212 473210 291240 488022
rect 291292 484152 291344 484158
rect 291292 484094 291344 484100
rect 291304 477426 291332 484094
rect 291488 478650 291516 488022
rect 291948 484158 291976 488022
rect 291936 484152 291988 484158
rect 291936 484094 291988 484100
rect 292580 480888 292632 480894
rect 292580 480830 292632 480836
rect 291476 478644 291528 478650
rect 291476 478586 291528 478592
rect 291292 477420 291344 477426
rect 291292 477362 291344 477368
rect 291200 473204 291252 473210
rect 291200 473146 291252 473152
rect 289820 470552 289872 470558
rect 289820 470494 289872 470500
rect 287060 470280 287112 470286
rect 287060 470222 287112 470228
rect 285772 470212 285824 470218
rect 285772 470154 285824 470160
rect 292592 467129 292620 480830
rect 292776 480214 292804 488022
rect 292868 488022 293158 488050
rect 293328 488022 293618 488050
rect 292764 480208 292816 480214
rect 292764 480150 292816 480156
rect 292868 476114 292896 488022
rect 293328 480894 293356 488022
rect 293988 487830 294016 488036
rect 294064 488022 294446 488050
rect 294616 488022 294906 488050
rect 293976 487824 294028 487830
rect 293976 487766 294028 487772
rect 293316 480888 293368 480894
rect 293316 480830 293368 480836
rect 293960 480888 294012 480894
rect 293960 480830 294012 480836
rect 292684 476086 292896 476114
rect 292684 467634 292712 476086
rect 292672 467628 292724 467634
rect 292672 467570 292724 467576
rect 292578 467120 292634 467129
rect 292578 467055 292634 467064
rect 285680 465588 285732 465594
rect 285680 465530 285732 465536
rect 293972 464438 294000 480830
rect 294064 468450 294092 488022
rect 294144 487824 294196 487830
rect 294144 487766 294196 487772
rect 294156 475561 294184 487766
rect 294616 480894 294644 488022
rect 294604 480888 294656 480894
rect 294604 480830 294656 480836
rect 294142 475552 294198 475561
rect 294142 475487 294198 475496
rect 295352 471578 295380 488036
rect 295444 488022 295826 488050
rect 295904 488022 296194 488050
rect 296272 488022 296654 488050
rect 296732 488022 297114 488050
rect 297192 488022 297574 488050
rect 297744 488022 298034 488050
rect 298112 488022 298402 488050
rect 298480 488022 298862 488050
rect 299338 488022 299428 488050
rect 295444 471850 295472 488022
rect 295524 480888 295576 480894
rect 295524 480830 295576 480836
rect 295536 471918 295564 480830
rect 295904 471986 295932 488022
rect 296272 480894 296300 488022
rect 296260 480888 296312 480894
rect 296260 480830 296312 480836
rect 295892 471980 295944 471986
rect 295892 471922 295944 471928
rect 295524 471912 295576 471918
rect 295524 471854 295576 471860
rect 295432 471844 295484 471850
rect 295432 471786 295484 471792
rect 296732 471714 296760 488022
rect 297192 477057 297220 488022
rect 297744 480078 297772 488022
rect 297732 480072 297784 480078
rect 297732 480014 297784 480020
rect 297178 477048 297234 477057
rect 297178 476983 297234 476992
rect 296720 471708 296772 471714
rect 296720 471650 296772 471656
rect 298112 471646 298140 488022
rect 298480 478514 298508 488022
rect 299400 482934 299428 488022
rect 299492 488022 299782 488050
rect 299388 482928 299440 482934
rect 299388 482870 299440 482876
rect 298468 478508 298520 478514
rect 298468 478450 298520 478456
rect 298100 471640 298152 471646
rect 298100 471582 298152 471588
rect 295340 471572 295392 471578
rect 295340 471514 295392 471520
rect 299492 471170 299520 488022
rect 316696 482225 316724 616830
rect 316788 552906 316816 635326
rect 316960 634024 317012 634030
rect 316960 633966 317012 633972
rect 316868 633480 316920 633486
rect 316868 633422 316920 633428
rect 316880 568410 316908 633422
rect 316868 568404 316920 568410
rect 316868 568346 316920 568352
rect 316972 568342 317000 633966
rect 317052 632256 317104 632262
rect 317052 632198 317104 632204
rect 316960 568336 317012 568342
rect 316960 568278 317012 568284
rect 317064 568274 317092 632198
rect 317144 579692 317196 579698
rect 317144 579634 317196 579640
rect 317052 568268 317104 568274
rect 317052 568210 317104 568216
rect 317156 566778 317184 579634
rect 317144 566772 317196 566778
rect 317144 566714 317196 566720
rect 318076 562562 318104 635530
rect 318168 569906 318196 638182
rect 320824 636880 320876 636886
rect 320824 636822 320876 636828
rect 319444 635452 319496 635458
rect 319444 635394 319496 635400
rect 318156 569900 318208 569906
rect 318156 569842 318208 569848
rect 318064 562556 318116 562562
rect 318064 562498 318116 562504
rect 319456 559638 319484 635394
rect 319628 632392 319680 632398
rect 319628 632334 319680 632340
rect 319536 632188 319588 632194
rect 319536 632130 319588 632136
rect 319548 567798 319576 632130
rect 319640 568138 319668 632334
rect 319628 568132 319680 568138
rect 319628 568074 319680 568080
rect 319536 567792 319588 567798
rect 319536 567734 319588 567740
rect 319444 559632 319496 559638
rect 319444 559574 319496 559580
rect 316776 552900 316828 552906
rect 316776 552842 316828 552848
rect 316960 552492 317012 552498
rect 316960 552434 317012 552440
rect 316868 552424 316920 552430
rect 316868 552366 316920 552372
rect 316776 550928 316828 550934
rect 316776 550870 316828 550876
rect 316788 518770 316816 550870
rect 316776 518764 316828 518770
rect 316776 518706 316828 518712
rect 316880 517342 316908 552366
rect 316972 517410 317000 552434
rect 317052 552288 317104 552294
rect 317052 552230 317104 552236
rect 317064 518838 317092 552230
rect 319444 552220 319496 552226
rect 319444 552162 319496 552168
rect 318064 550996 318116 551002
rect 318064 550938 318116 550944
rect 317144 550860 317196 550866
rect 317144 550802 317196 550808
rect 317156 518906 317184 550802
rect 317234 548040 317290 548049
rect 317234 547975 317290 547984
rect 317144 518900 317196 518906
rect 317144 518842 317196 518848
rect 317052 518832 317104 518838
rect 317052 518774 317104 518780
rect 316960 517404 317012 517410
rect 316960 517346 317012 517352
rect 316868 517336 316920 517342
rect 316868 517278 316920 517284
rect 317248 517274 317276 547975
rect 318076 520266 318104 550938
rect 319456 521558 319484 552162
rect 320836 550633 320864 636822
rect 355600 635792 355652 635798
rect 355600 635734 355652 635740
rect 322480 635724 322532 635730
rect 322480 635666 322532 635672
rect 346584 635724 346636 635730
rect 346584 635666 346636 635672
rect 322296 635656 322348 635662
rect 322296 635598 322348 635604
rect 321008 635112 321060 635118
rect 321008 635054 321060 635060
rect 320916 633548 320968 633554
rect 320916 633490 320968 633496
rect 320822 550624 320878 550633
rect 320822 550559 320878 550568
rect 320928 550225 320956 633490
rect 321020 554266 321048 635054
rect 322204 633616 322256 633622
rect 322204 633558 322256 633564
rect 321098 632224 321154 632233
rect 321098 632159 321154 632168
rect 321112 565146 321140 632159
rect 321558 627464 321614 627473
rect 321558 627399 321614 627408
rect 321572 626618 321600 627399
rect 321560 626612 321612 626618
rect 321560 626554 321612 626560
rect 321558 622704 321614 622713
rect 321558 622639 321614 622648
rect 321572 622470 321600 622639
rect 321560 622464 321612 622470
rect 321560 622406 321612 622412
rect 321558 617944 321614 617953
rect 321558 617879 321614 617888
rect 321572 616894 321600 617879
rect 321560 616888 321612 616894
rect 321560 616830 321612 616836
rect 321558 613184 321614 613193
rect 321558 613119 321614 613128
rect 321572 612814 321600 613119
rect 321560 612808 321612 612814
rect 321560 612750 321612 612756
rect 321558 608424 321614 608433
rect 321558 608359 321614 608368
rect 321572 607238 321600 608359
rect 321560 607232 321612 607238
rect 321560 607174 321612 607180
rect 321558 603664 321614 603673
rect 321558 603599 321614 603608
rect 321572 603158 321600 603599
rect 321560 603152 321612 603158
rect 321560 603094 321612 603100
rect 321558 598904 321614 598913
rect 321558 598839 321614 598848
rect 321572 597582 321600 598839
rect 321560 597576 321612 597582
rect 321560 597518 321612 597524
rect 321558 589384 321614 589393
rect 321558 589319 321560 589328
rect 321612 589319 321614 589328
rect 321560 589290 321612 589296
rect 321558 584624 321614 584633
rect 321558 584559 321614 584568
rect 321572 583778 321600 584559
rect 321560 583772 321612 583778
rect 321560 583714 321612 583720
rect 321558 579864 321614 579873
rect 321558 579799 321614 579808
rect 321572 579698 321600 579799
rect 321560 579692 321612 579698
rect 321560 579634 321612 579640
rect 321558 574424 321614 574433
rect 321558 574359 321614 574368
rect 321572 574122 321600 574359
rect 321560 574116 321612 574122
rect 321560 574058 321612 574064
rect 321560 569900 321612 569906
rect 321560 569842 321612 569848
rect 321572 569673 321600 569842
rect 321558 569664 321614 569673
rect 321558 569599 321614 569608
rect 321100 565140 321152 565146
rect 321100 565082 321152 565088
rect 321558 564904 321614 564913
rect 321558 564839 321614 564848
rect 321572 563718 321600 564839
rect 321560 563712 321612 563718
rect 321560 563654 321612 563660
rect 321558 560144 321614 560153
rect 321558 560079 321614 560088
rect 321572 558958 321600 560079
rect 321560 558952 321612 558958
rect 321560 558894 321612 558900
rect 321558 555384 321614 555393
rect 321558 555319 321614 555328
rect 321572 554810 321600 555319
rect 321560 554804 321612 554810
rect 321560 554746 321612 554752
rect 321008 554260 321060 554266
rect 321008 554202 321060 554208
rect 321008 551132 321060 551138
rect 321008 551074 321060 551080
rect 320914 550216 320970 550225
rect 320914 550151 320970 550160
rect 319536 549636 319588 549642
rect 319536 549578 319588 549584
rect 319444 521552 319496 521558
rect 319444 521494 319496 521500
rect 319548 521150 319576 549578
rect 319720 549568 319772 549574
rect 319720 549510 319772 549516
rect 319628 549500 319680 549506
rect 319628 549442 319680 549448
rect 319640 521422 319668 549442
rect 319628 521416 319680 521422
rect 319628 521358 319680 521364
rect 319536 521144 319588 521150
rect 319536 521086 319588 521092
rect 319732 520742 319760 549510
rect 319812 548820 319864 548826
rect 319812 548762 319864 548768
rect 319824 521490 319852 548762
rect 320824 539640 320876 539646
rect 320824 539582 320876 539588
rect 319812 521484 319864 521490
rect 319812 521426 319864 521432
rect 319720 520736 319772 520742
rect 319720 520678 319772 520684
rect 318064 520260 318116 520266
rect 318064 520202 318116 520208
rect 317236 517268 317288 517274
rect 317236 517210 317288 517216
rect 320836 489190 320864 539582
rect 321020 519654 321048 551074
rect 322216 550089 322244 633558
rect 322308 562698 322336 635598
rect 322388 634908 322440 634914
rect 322388 634850 322440 634856
rect 322400 563922 322428 634850
rect 322492 565214 322520 635666
rect 323952 635520 324004 635526
rect 323952 635462 324004 635468
rect 323860 634976 323912 634982
rect 323860 634918 323912 634924
rect 323768 634840 323820 634846
rect 323768 634782 323820 634788
rect 323676 634364 323728 634370
rect 323676 634306 323728 634312
rect 322572 634296 322624 634302
rect 322572 634238 322624 634244
rect 322584 568070 322612 634238
rect 322664 634160 322716 634166
rect 322664 634102 322716 634108
rect 322676 596834 322704 634102
rect 323584 632460 323636 632466
rect 323584 632402 323636 632408
rect 322664 596828 322716 596834
rect 322664 596770 322716 596776
rect 322572 568064 322624 568070
rect 322572 568006 322624 568012
rect 322480 565208 322532 565214
rect 322480 565150 322532 565156
rect 322388 563916 322440 563922
rect 322388 563858 322440 563864
rect 322296 562692 322348 562698
rect 322296 562634 322348 562640
rect 322388 552152 322440 552158
rect 322388 552094 322440 552100
rect 322296 550724 322348 550730
rect 322296 550666 322348 550672
rect 322202 550080 322258 550089
rect 322202 550015 322258 550024
rect 321098 549400 321154 549409
rect 321098 549335 321154 549344
rect 321112 522646 321140 549335
rect 321836 548684 321888 548690
rect 321836 548626 321888 548632
rect 321848 545873 321876 548626
rect 322204 548548 322256 548554
rect 322204 548490 322256 548496
rect 321834 545864 321890 545873
rect 321834 545799 321890 545808
rect 321560 542360 321612 542366
rect 321560 542302 321612 542308
rect 321572 541113 321600 542302
rect 321558 541104 321614 541113
rect 321558 541039 321614 541048
rect 321560 536784 321612 536790
rect 321560 536726 321612 536732
rect 321572 536353 321600 536726
rect 321558 536344 321614 536353
rect 321558 536279 321614 536288
rect 322216 531593 322244 548490
rect 322202 531584 322258 531593
rect 322202 531519 322258 531528
rect 321560 527128 321612 527134
rect 321560 527070 321612 527076
rect 321572 526833 321600 527070
rect 321558 526824 321614 526833
rect 321558 526759 321614 526768
rect 321100 522640 321152 522646
rect 321100 522582 321152 522588
rect 322308 519994 322336 550666
rect 322400 521082 322428 552094
rect 322572 552084 322624 552090
rect 322572 552026 322624 552032
rect 322480 550792 322532 550798
rect 322480 550734 322532 550740
rect 322388 521076 322440 521082
rect 322388 521018 322440 521024
rect 322296 519988 322348 519994
rect 322296 519930 322348 519936
rect 322492 519722 322520 550734
rect 322584 521014 322612 552026
rect 322756 550180 322808 550186
rect 322756 550122 322808 550128
rect 322664 549432 322716 549438
rect 322664 549374 322716 549380
rect 322572 521008 322624 521014
rect 322572 520950 322624 520956
rect 322676 520946 322704 549374
rect 322768 522578 322796 550122
rect 322756 522572 322808 522578
rect 322756 522514 322808 522520
rect 323596 521626 323624 632402
rect 323688 549953 323716 634306
rect 323780 556986 323808 634782
rect 323872 558278 323900 634918
rect 323964 561202 323992 635462
rect 342260 635384 342312 635390
rect 342260 635326 342312 635332
rect 324872 635316 324924 635322
rect 324872 635258 324924 635264
rect 324778 634944 324834 634953
rect 324778 634879 324834 634888
rect 324228 634092 324280 634098
rect 324228 634034 324280 634040
rect 324240 594153 324268 634034
rect 324226 594144 324282 594153
rect 324226 594079 324282 594088
rect 324792 562630 324820 634879
rect 324780 562624 324832 562630
rect 324780 562566 324832 562572
rect 323952 561196 324004 561202
rect 323952 561138 324004 561144
rect 323860 558272 323912 558278
rect 323860 558214 323912 558220
rect 323768 556980 323820 556986
rect 323768 556922 323820 556928
rect 324884 552838 324912 635258
rect 337568 634908 337620 634914
rect 337568 634850 337620 634856
rect 328644 634840 328696 634846
rect 328644 634782 328696 634788
rect 328656 633026 328684 634782
rect 337580 633026 337608 634850
rect 342272 633026 342300 635326
rect 346596 633026 346624 635666
rect 353300 635248 353352 635254
rect 353300 635190 353352 635196
rect 328656 632998 328900 633026
rect 337580 632998 337916 633026
rect 342272 632998 342424 633026
rect 346596 632998 346932 633026
rect 353312 632874 353340 635190
rect 355612 633026 355640 635734
rect 392308 635588 392360 635594
rect 392308 635530 392360 635536
rect 369124 635520 369176 635526
rect 369124 635462 369176 635468
rect 364616 635452 364668 635458
rect 364616 635394 364668 635400
rect 361396 635384 361448 635390
rect 361396 635326 361448 635332
rect 360200 634228 360252 634234
rect 360200 634170 360252 634176
rect 360212 633026 360240 634170
rect 355612 632998 355948 633026
rect 360212 632998 360456 633026
rect 353300 632868 353352 632874
rect 353300 632810 353352 632816
rect 361408 632806 361436 635326
rect 364628 633026 364656 635394
rect 369136 633026 369164 635462
rect 378140 635316 378192 635322
rect 378140 635258 378192 635264
rect 374000 635180 374052 635186
rect 374000 635122 374052 635128
rect 374012 633026 374040 635122
rect 364628 632998 364964 633026
rect 369136 632998 369472 633026
rect 373980 632998 374040 633026
rect 378152 633026 378180 635258
rect 387800 635112 387852 635118
rect 387800 635054 387852 635060
rect 383660 635044 383712 635050
rect 383660 634986 383712 634992
rect 383672 633026 383700 634986
rect 378152 632998 378488 633026
rect 383640 632998 383700 633026
rect 387812 633026 387840 635054
rect 391940 634840 391992 634846
rect 391940 634782 391992 634788
rect 387812 632998 388148 633026
rect 361396 632800 361448 632806
rect 361396 632742 361448 632748
rect 391952 632738 391980 634782
rect 392320 633026 392348 635530
rect 401600 634976 401652 634982
rect 401600 634918 401652 634924
rect 396816 633820 396868 633826
rect 396816 633762 396868 633768
rect 396828 633026 396856 633762
rect 401612 633298 401640 634918
rect 401612 633270 401686 633298
rect 392320 632998 392656 633026
rect 396828 632998 397164 633026
rect 401658 633012 401686 633270
rect 405752 633026 405780 640970
rect 428280 638240 428332 638246
rect 428280 638182 428332 638188
rect 414848 635384 414900 635390
rect 414848 635326 414900 635332
rect 410340 635248 410392 635254
rect 410340 635190 410392 635196
rect 410352 633026 410380 635190
rect 414860 633026 414888 635326
rect 423862 634944 423918 634953
rect 423862 634879 423918 634888
rect 420000 634840 420052 634846
rect 420000 634782 420052 634788
rect 420012 633026 420040 634782
rect 405752 632998 406180 633026
rect 410352 632998 410688 633026
rect 414860 632998 415196 633026
rect 419704 632998 420040 633026
rect 423876 633026 423904 634879
rect 428292 633026 428320 638182
rect 432880 635656 432932 635662
rect 432880 635598 432932 635604
rect 432892 633026 432920 635598
rect 423876 632998 424212 633026
rect 428292 632998 428720 633026
rect 432892 632998 433228 633026
rect 391940 632732 391992 632738
rect 391940 632674 391992 632680
rect 333058 632632 333114 632641
rect 333114 632590 333408 632618
rect 333058 632567 333114 632576
rect 351090 632496 351146 632505
rect 351146 632454 351440 632482
rect 351090 632431 351146 632440
rect 433340 632324 433392 632330
rect 433340 632266 433392 632272
rect 433352 619177 433380 632266
rect 433338 619168 433394 619177
rect 433338 619103 433394 619112
rect 433338 589520 433394 589529
rect 433338 589455 433394 589464
rect 324872 552832 324924 552838
rect 324872 552774 324924 552780
rect 323768 551064 323820 551070
rect 323768 551006 323820 551012
rect 323674 549944 323730 549953
rect 323674 549879 323730 549888
rect 323676 548344 323728 548350
rect 323676 548286 323728 548292
rect 323584 521620 323636 521626
rect 323584 521562 323636 521568
rect 322664 520940 322716 520946
rect 322664 520882 322716 520888
rect 323688 520334 323716 548286
rect 323676 520328 323728 520334
rect 323676 520270 323728 520276
rect 323780 519858 323808 551006
rect 324872 550656 324924 550662
rect 324872 550598 324924 550604
rect 323952 550112 324004 550118
rect 323952 550054 324004 550060
rect 323860 548072 323912 548078
rect 323860 548014 323912 548020
rect 323872 520198 323900 548014
rect 323964 522510 323992 550054
rect 324780 548412 324832 548418
rect 324780 548354 324832 548360
rect 324688 548140 324740 548146
rect 324688 548082 324740 548088
rect 324700 528554 324728 548082
rect 324516 528526 324728 528554
rect 323952 522504 324004 522510
rect 323952 522446 324004 522452
rect 323860 520192 323912 520198
rect 323860 520134 323912 520140
rect 323768 519852 323820 519858
rect 323768 519794 323820 519800
rect 322480 519716 322532 519722
rect 322480 519658 322532 519664
rect 321008 519648 321060 519654
rect 321008 519590 321060 519596
rect 324516 519586 324544 528526
rect 324792 524362 324820 548354
rect 324608 524334 324820 524362
rect 324608 520130 324636 524334
rect 324884 522442 324912 550598
rect 324872 522436 324924 522442
rect 324872 522378 324924 522384
rect 325148 522436 325200 522442
rect 325148 522378 325200 522384
rect 324700 522294 325036 522322
rect 324700 520266 324728 522294
rect 324688 520260 324740 520266
rect 324688 520202 324740 520208
rect 324596 520124 324648 520130
rect 324596 520066 324648 520072
rect 324504 519580 324556 519586
rect 324504 519522 324556 519528
rect 325160 519382 325188 522378
rect 329544 522022 329788 522050
rect 334052 522022 334112 522050
rect 329760 520033 329788 522022
rect 334084 520130 334112 522022
rect 338224 522022 338560 522050
rect 342732 522022 343068 522050
rect 347240 522022 347576 522050
rect 351932 522022 352084 522050
rect 356256 522022 356592 522050
rect 360212 522022 361100 522050
rect 365272 522022 365608 522050
rect 369872 522022 370116 522050
rect 374288 522022 374624 522050
rect 379532 522022 379776 522050
rect 383672 522022 384284 522050
rect 388456 522022 388792 522050
rect 393300 522022 393360 522050
rect 338224 520198 338252 522022
rect 342732 521626 342760 522022
rect 342720 521620 342772 521626
rect 342720 521562 342772 521568
rect 347240 520266 347268 522022
rect 347228 520260 347280 520266
rect 347228 520202 347280 520208
rect 338212 520192 338264 520198
rect 338212 520134 338264 520140
rect 334072 520124 334124 520130
rect 334072 520066 334124 520072
rect 329746 520024 329802 520033
rect 329746 519959 329802 519968
rect 351932 519586 351960 522022
rect 356256 520810 356284 522022
rect 356244 520804 356296 520810
rect 356244 520746 356296 520752
rect 351920 519580 351972 519586
rect 351920 519522 351972 519528
rect 325148 519376 325200 519382
rect 325148 519318 325200 519324
rect 320824 489184 320876 489190
rect 320824 489126 320876 489132
rect 360212 488102 360240 522022
rect 365272 519790 365300 522022
rect 365260 519784 365312 519790
rect 365260 519726 365312 519732
rect 369872 519654 369900 522022
rect 374288 520878 374316 522022
rect 374276 520872 374328 520878
rect 374276 520814 374328 520820
rect 379532 519722 379560 522022
rect 379520 519716 379572 519722
rect 379520 519658 379572 519664
rect 369860 519648 369912 519654
rect 369860 519590 369912 519596
rect 360200 488096 360252 488102
rect 360200 488038 360252 488044
rect 356612 486532 356664 486538
rect 356612 486474 356664 486480
rect 316682 482216 316738 482225
rect 316682 482151 316738 482160
rect 299480 471164 299532 471170
rect 299480 471106 299532 471112
rect 294052 468444 294104 468450
rect 294052 468386 294104 468392
rect 339408 466608 339460 466614
rect 338486 466576 338542 466585
rect 339408 466550 339460 466556
rect 339774 466576 339830 466585
rect 338486 466511 338542 466520
rect 338500 466478 338528 466511
rect 339420 466478 339448 466550
rect 339774 466511 339776 466520
rect 339828 466511 339830 466520
rect 350998 466576 351054 466585
rect 350998 466511 351054 466520
rect 339776 466482 339828 466488
rect 351012 466478 351040 466511
rect 338488 466472 338540 466478
rect 338488 466414 338540 466420
rect 339408 466472 339460 466478
rect 339408 466414 339460 466420
rect 351000 466472 351052 466478
rect 351000 466414 351052 466420
rect 293960 464432 294012 464438
rect 293960 464374 294012 464380
rect 271880 464364 271932 464370
rect 271880 464306 271932 464312
rect 256056 380996 256108 381002
rect 256056 380938 256108 380944
rect 256068 380769 256096 380938
rect 235998 380760 236054 380769
rect 235998 380695 236054 380704
rect 237102 380760 237158 380769
rect 237102 380695 237158 380704
rect 243082 380760 243138 380769
rect 243082 380695 243138 380704
rect 245382 380760 245438 380769
rect 245382 380695 245438 380704
rect 256054 380760 256110 380769
rect 256054 380695 256110 380704
rect 269762 380760 269818 380769
rect 269762 380695 269818 380704
rect 236012 379982 236040 380695
rect 236000 379976 236052 379982
rect 236000 379918 236052 379924
rect 237116 379846 237144 380695
rect 240048 379976 240100 379982
rect 240048 379918 240100 379924
rect 237104 379840 237156 379846
rect 237104 379782 237156 379788
rect 237380 379840 237432 379846
rect 237380 379782 237432 379788
rect 220820 379772 220872 379778
rect 220820 379714 220872 379720
rect 220832 379658 220860 379714
rect 221004 379704 221056 379710
rect 220832 379652 221004 379658
rect 220832 379646 221056 379652
rect 220832 379630 221044 379646
rect 220268 379364 220320 379370
rect 220268 379306 220320 379312
rect 220280 378350 220308 379306
rect 220728 379228 220780 379234
rect 220728 379170 220780 379176
rect 220740 378690 220768 379170
rect 220912 379160 220964 379166
rect 220912 379102 220964 379108
rect 220820 378888 220872 378894
rect 220820 378830 220872 378836
rect 220728 378684 220780 378690
rect 220728 378626 220780 378632
rect 220268 378344 220320 378350
rect 220268 378286 220320 378292
rect 220832 358562 220860 378830
rect 220924 378350 220952 379102
rect 221188 379092 221240 379098
rect 221188 379034 221240 379040
rect 222016 379092 222068 379098
rect 222016 379034 222068 379040
rect 221004 379024 221056 379030
rect 221004 378966 221056 378972
rect 220912 378344 220964 378350
rect 220912 378286 220964 378292
rect 220820 358556 220872 358562
rect 220820 358498 220872 358504
rect 220924 357610 220952 378286
rect 221016 358698 221044 378966
rect 221094 378448 221150 378457
rect 221094 378383 221150 378392
rect 221004 358692 221056 358698
rect 221004 358634 221056 358640
rect 221108 358222 221136 378383
rect 221200 358766 221228 379034
rect 221280 378616 221332 378622
rect 221280 378558 221332 378564
rect 221188 358760 221240 358766
rect 221188 358702 221240 358708
rect 221292 358290 221320 378558
rect 222028 378486 222056 379034
rect 222108 378888 222160 378894
rect 222108 378830 222160 378836
rect 222016 378480 222068 378486
rect 222016 378422 222068 378428
rect 222120 378418 222148 378830
rect 222108 378412 222160 378418
rect 222108 378354 222160 378360
rect 237392 377534 237420 379782
rect 237380 377528 237432 377534
rect 237380 377470 237432 377476
rect 240060 375834 240088 379918
rect 243096 379914 243124 380695
rect 243084 379908 243136 379914
rect 243084 379850 243136 379856
rect 245396 378826 245424 380695
rect 254490 380624 254546 380633
rect 254490 380559 254546 380568
rect 255870 380624 255926 380633
rect 255870 380559 255926 380568
rect 256974 380624 257030 380633
rect 256974 380559 257030 380568
rect 259458 380624 259514 380633
rect 259458 380559 259514 380568
rect 265254 380624 265310 380633
rect 265254 380559 265310 380568
rect 254504 379778 254532 380559
rect 254492 379772 254544 379778
rect 254492 379714 254544 379720
rect 255884 379710 255912 380559
rect 255872 379704 255924 379710
rect 255872 379646 255924 379652
rect 256988 379642 257016 380559
rect 259472 379982 259500 380559
rect 262864 380384 262916 380390
rect 262864 380326 262916 380332
rect 259460 379976 259512 379982
rect 259460 379918 259512 379924
rect 256976 379636 257028 379642
rect 256976 379578 257028 379584
rect 258080 379568 258132 379574
rect 258080 379510 258132 379516
rect 258092 379409 258120 379510
rect 246026 379400 246082 379409
rect 246026 379335 246082 379344
rect 247498 379400 247554 379409
rect 247498 379335 247554 379344
rect 248602 379400 248658 379409
rect 248602 379335 248658 379344
rect 250074 379400 250130 379409
rect 250074 379335 250130 379344
rect 251178 379400 251234 379409
rect 251178 379335 251234 379344
rect 252282 379400 252338 379409
rect 252282 379335 252338 379344
rect 253386 379400 253442 379409
rect 253386 379335 253442 379344
rect 258078 379400 258134 379409
rect 258078 379335 258134 379344
rect 261666 379400 261722 379409
rect 261666 379335 261722 379344
rect 245384 378820 245436 378826
rect 245384 378762 245436 378768
rect 246040 378758 246068 379335
rect 246028 378752 246080 378758
rect 246028 378694 246080 378700
rect 247512 378690 247540 379335
rect 248234 378856 248290 378865
rect 248234 378791 248290 378800
rect 247500 378684 247552 378690
rect 247500 378626 247552 378632
rect 244278 378312 244334 378321
rect 244278 378247 244334 378256
rect 240048 375828 240100 375834
rect 240048 375770 240100 375776
rect 244292 375018 244320 378247
rect 248248 376174 248276 378791
rect 248616 378554 248644 379335
rect 250088 378622 250116 379335
rect 250076 378616 250128 378622
rect 250076 378558 250128 378564
rect 248604 378548 248656 378554
rect 248604 378490 248656 378496
rect 251192 378486 251220 379335
rect 251180 378480 251232 378486
rect 251180 378422 251232 378428
rect 252296 378418 252324 379335
rect 253400 379302 253428 379335
rect 253388 379296 253440 379302
rect 253388 379238 253440 379244
rect 252374 378856 252430 378865
rect 252374 378791 252430 378800
rect 252388 378457 252416 378791
rect 253570 378584 253626 378593
rect 253570 378519 253626 378528
rect 258354 378584 258410 378593
rect 258354 378519 258410 378528
rect 260930 378584 260986 378593
rect 260930 378519 260986 378528
rect 252374 378448 252430 378457
rect 252284 378412 252336 378418
rect 252374 378383 252430 378392
rect 252284 378354 252336 378360
rect 250626 378312 250682 378321
rect 250626 378247 250682 378256
rect 248236 376168 248288 376174
rect 248236 376110 248288 376116
rect 250640 375902 250668 378247
rect 253584 375970 253612 378519
rect 258368 376038 258396 378519
rect 260944 376106 260972 378519
rect 260932 376100 260984 376106
rect 260932 376042 260984 376048
rect 258356 376032 258408 376038
rect 258356 375974 258408 375980
rect 253572 375964 253624 375970
rect 253572 375906 253624 375912
rect 250628 375896 250680 375902
rect 250628 375838 250680 375844
rect 261680 375154 261708 379335
rect 262876 378457 262904 380326
rect 265268 379846 265296 380559
rect 269776 380390 269804 380695
rect 270958 380624 271014 380633
rect 270958 380559 271014 380568
rect 269764 380384 269816 380390
rect 269764 380326 269816 380332
rect 265256 379840 265308 379846
rect 265256 379782 265308 379788
rect 268660 379432 268712 379438
rect 268658 379400 268660 379409
rect 268712 379400 268714 379409
rect 268658 379335 268714 379344
rect 263598 378584 263654 378593
rect 263598 378519 263654 378528
rect 265898 378584 265954 378593
rect 265898 378519 265954 378528
rect 268106 378584 268162 378593
rect 268106 378519 268162 378528
rect 262862 378448 262918 378457
rect 262862 378383 262918 378392
rect 262770 378312 262826 378321
rect 262770 378247 262826 378256
rect 262784 375222 262812 378247
rect 263612 376310 263640 378519
rect 265912 376378 265940 378519
rect 266358 378312 266414 378321
rect 266358 378247 266414 378256
rect 267554 378312 267610 378321
rect 267554 378247 267610 378256
rect 265900 376372 265952 376378
rect 265900 376314 265952 376320
rect 263600 376304 263652 376310
rect 263600 376246 263652 376252
rect 262772 375216 262824 375222
rect 262772 375158 262824 375164
rect 261668 375148 261720 375154
rect 261668 375090 261720 375096
rect 244280 375012 244332 375018
rect 244280 374954 244332 374960
rect 266372 374678 266400 378247
rect 267568 375290 267596 378247
rect 268120 376446 268148 378519
rect 268108 376440 268160 376446
rect 268108 376382 268160 376388
rect 270972 376242 271000 380559
rect 274640 380452 274692 380458
rect 274640 380394 274692 380400
rect 274652 379506 274680 380394
rect 293960 380316 294012 380322
rect 293960 380258 294012 380264
rect 273260 379500 273312 379506
rect 273260 379442 273312 379448
rect 274640 379500 274692 379506
rect 274640 379442 274692 379448
rect 273272 379409 273300 379442
rect 271050 379400 271106 379409
rect 271050 379335 271052 379344
rect 271104 379335 271106 379344
rect 272062 379400 272118 379409
rect 272062 379335 272118 379344
rect 273258 379400 273314 379409
rect 273258 379335 273314 379344
rect 274178 379400 274234 379409
rect 274178 379335 274234 379344
rect 275650 379400 275706 379409
rect 275650 379335 275706 379344
rect 276018 379400 276074 379409
rect 276018 379335 276074 379344
rect 276938 379400 276994 379409
rect 276938 379335 276994 379344
rect 285954 379400 286010 379409
rect 285954 379335 286010 379344
rect 287702 379400 287758 379409
rect 287702 379335 287758 379344
rect 290922 379400 290978 379409
rect 290922 379335 290978 379344
rect 292670 379400 292726 379409
rect 292670 379335 292726 379344
rect 271052 379306 271104 379312
rect 272076 378282 272104 379335
rect 273442 378584 273498 378593
rect 273442 378519 273498 378528
rect 272064 378276 272116 378282
rect 272064 378218 272116 378224
rect 273456 376582 273484 378519
rect 274192 378350 274220 379335
rect 274180 378344 274232 378350
rect 274180 378286 274232 378292
rect 274272 378344 274324 378350
rect 274272 378286 274324 378292
rect 274284 377330 274312 378286
rect 275664 378214 275692 379335
rect 274640 378208 274692 378214
rect 274638 378176 274640 378185
rect 275652 378208 275704 378214
rect 274692 378176 274694 378185
rect 275652 378150 275704 378156
rect 274638 378111 274694 378120
rect 274272 377324 274324 377330
rect 274272 377266 274324 377272
rect 273444 376576 273496 376582
rect 273444 376518 273496 376524
rect 276032 376514 276060 379335
rect 276952 378894 276980 379335
rect 277858 379264 277914 379273
rect 277858 379199 277914 379208
rect 278042 379264 278098 379273
rect 278042 379199 278098 379208
rect 279146 379264 279202 379273
rect 279146 379199 279202 379208
rect 280710 379264 280766 379273
rect 280710 379199 280766 379208
rect 283010 379264 283066 379273
rect 283010 379199 283066 379208
rect 276940 378888 276992 378894
rect 276940 378830 276992 378836
rect 277872 378282 277900 379199
rect 277860 378276 277912 378282
rect 277860 378218 277912 378224
rect 278056 377398 278084 379199
rect 278044 377392 278096 377398
rect 278044 377334 278096 377340
rect 276020 376508 276072 376514
rect 276020 376450 276072 376456
rect 270960 376236 271012 376242
rect 270960 376178 271012 376184
rect 267556 375284 267608 375290
rect 267556 375226 267608 375232
rect 279160 375086 279188 379199
rect 280724 377466 280752 379199
rect 280712 377460 280764 377466
rect 280712 377402 280764 377408
rect 283024 376718 283052 379199
rect 285968 377602 285996 379335
rect 287716 377670 287744 379335
rect 290936 377738 290964 379335
rect 292684 377806 292712 379335
rect 293972 379302 294000 380258
rect 301504 380248 301556 380254
rect 301504 380190 301556 380196
rect 295890 379400 295946 379409
rect 295890 379335 295946 379344
rect 298466 379400 298522 379409
rect 298466 379335 298522 379344
rect 300858 379400 300914 379409
rect 301516 379370 301544 380190
rect 309048 380180 309100 380186
rect 309048 380122 309100 380128
rect 309060 379438 309088 380122
rect 356624 379506 356652 486474
rect 383672 486470 383700 522022
rect 388456 519926 388484 522022
rect 393332 520062 393360 522022
rect 397472 522022 397808 522050
rect 401980 522022 402316 522050
rect 406488 522022 406824 522050
rect 411332 522022 411392 522050
rect 393320 520056 393372 520062
rect 393320 519998 393372 520004
rect 388444 519920 388496 519926
rect 388444 519862 388496 519868
rect 397472 516769 397500 522022
rect 401980 519858 402008 522022
rect 406488 519994 406516 522022
rect 406476 519988 406528 519994
rect 406476 519930 406528 519936
rect 401968 519852 402020 519858
rect 401968 519794 402020 519800
rect 411364 519450 411392 522022
rect 415504 522022 415840 522050
rect 420012 522022 420348 522050
rect 424520 522022 424856 522050
rect 429212 522022 429364 522050
rect 415504 519518 415532 522022
rect 420012 521218 420040 522022
rect 420000 521212 420052 521218
rect 420000 521154 420052 521160
rect 415492 519512 415544 519518
rect 415492 519454 415544 519460
rect 411352 519444 411404 519450
rect 411352 519386 411404 519392
rect 424520 519382 424548 522022
rect 429212 520169 429240 522022
rect 433352 520946 433380 589455
rect 433430 574560 433486 574569
rect 433430 574495 433486 574504
rect 433444 521150 433472 574495
rect 433522 560416 433578 560425
rect 433522 560351 433578 560360
rect 433536 523002 433564 560351
rect 433614 546408 433670 546417
rect 433614 546343 433670 546352
rect 433628 538214 433656 546343
rect 433628 538186 433748 538214
rect 433536 522974 433656 523002
rect 433524 522708 433576 522714
rect 433524 522650 433576 522656
rect 433536 522617 433564 522650
rect 433522 522608 433578 522617
rect 433522 522543 433578 522552
rect 433432 521144 433484 521150
rect 433432 521086 433484 521092
rect 433628 521014 433656 522974
rect 433720 521082 433748 538186
rect 433708 521076 433760 521082
rect 433708 521018 433760 521024
rect 433616 521008 433668 521014
rect 433616 520950 433668 520956
rect 433340 520940 433392 520946
rect 433340 520882 433392 520888
rect 429198 520160 429254 520169
rect 429198 520095 429254 520104
rect 434732 520033 434760 700402
rect 434904 700392 434956 700398
rect 434904 700334 434956 700340
rect 434812 639600 434864 639606
rect 434812 639542 434864 639548
rect 434824 532273 434852 639542
rect 434916 628153 434944 700334
rect 457444 634840 457496 634846
rect 457444 634782 457496 634788
rect 436192 634364 436244 634370
rect 436192 634306 436244 634312
rect 436100 634296 436152 634302
rect 436100 634238 436152 634244
rect 434902 628144 434958 628153
rect 434902 628079 434958 628088
rect 436112 609113 436140 634238
rect 436204 613873 436232 634306
rect 456800 633956 456852 633962
rect 456800 633898 456852 633904
rect 436284 632392 436336 632398
rect 436284 632334 436336 632340
rect 436296 623393 436324 632334
rect 456812 627745 456840 633898
rect 456798 627736 456854 627745
rect 456798 627671 456854 627680
rect 436282 623384 436338 623393
rect 436282 623319 436338 623328
rect 436190 613864 436246 613873
rect 436190 613799 436246 613808
rect 436098 609104 436154 609113
rect 436098 609039 436154 609048
rect 436098 604344 436154 604353
rect 436098 604279 436154 604288
rect 434902 585304 434958 585313
rect 434902 585239 434958 585248
rect 434810 532264 434866 532273
rect 434810 532199 434866 532208
rect 434718 520024 434774 520033
rect 434718 519959 434774 519968
rect 424508 519376 424560 519382
rect 424508 519318 424560 519324
rect 397458 516760 397514 516769
rect 397458 516695 397514 516704
rect 383660 486464 383712 486470
rect 383660 486406 383712 486412
rect 356704 485580 356756 485586
rect 356704 485522 356756 485528
rect 323308 379500 323360 379506
rect 323308 379442 323360 379448
rect 325976 379500 326028 379506
rect 325976 379442 326028 379448
rect 356612 379500 356664 379506
rect 356612 379442 356664 379448
rect 309048 379432 309100 379438
rect 302790 379400 302846 379409
rect 300858 379335 300914 379344
rect 301504 379364 301556 379370
rect 293960 379296 294012 379302
rect 293960 379238 294012 379244
rect 295904 377874 295932 379335
rect 298480 378010 298508 379335
rect 300872 378078 300900 379335
rect 302790 379335 302846 379344
rect 305826 379400 305882 379409
rect 315764 379432 315816 379438
rect 309048 379374 309100 379380
rect 310978 379400 311034 379409
rect 305826 379335 305882 379344
rect 310978 379335 311034 379344
rect 313370 379400 313426 379409
rect 313370 379335 313372 379344
rect 301504 379306 301556 379312
rect 302804 378350 302832 379335
rect 302792 378344 302844 378350
rect 302792 378286 302844 378292
rect 300860 378072 300912 378078
rect 300860 378014 300912 378020
rect 298468 378004 298520 378010
rect 298468 377946 298520 377952
rect 305840 377942 305868 379335
rect 310992 379302 311020 379335
rect 313424 379335 313426 379344
rect 315762 379400 315764 379409
rect 323320 379409 323348 379442
rect 325988 379409 326016 379442
rect 315816 379400 315818 379409
rect 315762 379335 315818 379344
rect 317418 379400 317474 379409
rect 317418 379335 317474 379344
rect 323306 379400 323362 379409
rect 323306 379335 323362 379344
rect 325974 379400 326030 379409
rect 325974 379335 326030 379344
rect 343454 379400 343510 379409
rect 343454 379335 343510 379344
rect 313372 379306 313424 379312
rect 310980 379296 311032 379302
rect 310980 379238 311032 379244
rect 317432 378146 317460 379335
rect 320914 378584 320970 378593
rect 320914 378519 320970 378528
rect 317420 378140 317472 378146
rect 317420 378082 317472 378088
rect 305828 377936 305880 377942
rect 305828 377878 305880 377884
rect 295892 377868 295944 377874
rect 295892 377810 295944 377816
rect 292672 377800 292724 377806
rect 292672 377742 292724 377748
rect 290924 377732 290976 377738
rect 290924 377674 290976 377680
rect 287704 377664 287756 377670
rect 287704 377606 287756 377612
rect 285956 377596 286008 377602
rect 285956 377538 286008 377544
rect 283012 376712 283064 376718
rect 283012 376654 283064 376660
rect 320928 376650 320956 378519
rect 343178 378448 343234 378457
rect 343468 378418 343496 379335
rect 343178 378383 343234 378392
rect 343456 378412 343508 378418
rect 343192 378350 343220 378383
rect 343456 378354 343508 378360
rect 342260 378344 342312 378350
rect 342260 378286 342312 378292
rect 343180 378344 343232 378350
rect 343180 378286 343232 378292
rect 320916 376644 320968 376650
rect 320916 376586 320968 376592
rect 279148 375080 279200 375086
rect 279148 375022 279200 375028
rect 342272 374950 342300 378286
rect 356612 378208 356664 378214
rect 356612 378150 356664 378156
rect 342260 374944 342312 374950
rect 342260 374886 342312 374892
rect 266360 374672 266412 374678
rect 266360 374614 266412 374620
rect 339868 359576 339920 359582
rect 339868 359518 339920 359524
rect 339880 358873 339908 359518
rect 351736 359508 351788 359514
rect 351736 359450 351788 359456
rect 342260 358896 342312 358902
rect 338486 358864 338542 358873
rect 338486 358799 338488 358808
rect 338540 358799 338542 358808
rect 339866 358864 339922 358873
rect 351748 358873 351776 359450
rect 342260 358838 342312 358844
rect 351734 358864 351790 358873
rect 339866 358799 339922 358808
rect 338488 358770 338540 358776
rect 221280 358284 221332 358290
rect 221280 358226 221332 358232
rect 221096 358216 221148 358222
rect 221096 358158 221148 358164
rect 342272 358086 342300 358838
rect 351734 358799 351790 358808
rect 342260 358080 342312 358086
rect 342260 358022 342312 358028
rect 220912 357604 220964 357610
rect 220912 357546 220964 357552
rect 273168 273964 273220 273970
rect 273168 273906 273220 273912
rect 273180 273873 273208 273906
rect 273166 273864 273222 273873
rect 273166 273799 273222 273808
rect 266358 273592 266414 273601
rect 220820 273556 220872 273562
rect 266358 273527 266360 273536
rect 220820 273498 220872 273504
rect 266412 273527 266414 273536
rect 269762 273592 269818 273601
rect 269762 273527 269818 273536
rect 271142 273592 271198 273601
rect 271142 273527 271198 273536
rect 283470 273592 283526 273601
rect 283470 273527 283526 273536
rect 266360 273498 266412 273504
rect 220268 270428 220320 270434
rect 220268 270370 220320 270376
rect 220280 269346 220308 270370
rect 220636 270224 220688 270230
rect 220636 270166 220688 270172
rect 220268 269340 220320 269346
rect 220268 269282 220320 269288
rect 220648 269278 220676 270166
rect 220728 270156 220780 270162
rect 220728 270098 220780 270104
rect 220740 269618 220768 270098
rect 220728 269612 220780 269618
rect 220728 269554 220780 269560
rect 220636 269272 220688 269278
rect 220636 269214 220688 269220
rect 220832 252550 220860 273498
rect 269776 273494 269804 273527
rect 269764 273488 269816 273494
rect 269764 273430 269816 273436
rect 271156 273426 271184 273527
rect 273258 273456 273314 273465
rect 271144 273420 271196 273426
rect 273258 273391 273314 273400
rect 271144 273362 271196 273368
rect 273272 273358 273300 273391
rect 273260 273352 273312 273358
rect 273260 273294 273312 273300
rect 283484 273290 283512 273527
rect 283472 273284 283524 273290
rect 283472 273226 283524 273232
rect 285956 273148 286008 273154
rect 285956 273090 286008 273096
rect 285968 272921 285996 273090
rect 288164 273080 288216 273086
rect 288164 273022 288216 273028
rect 298466 273048 298522 273057
rect 288176 272921 288204 273022
rect 298466 272983 298468 272992
rect 298520 272983 298522 272992
rect 298468 272954 298520 272960
rect 295892 272944 295944 272950
rect 285954 272912 286010 272921
rect 285954 272847 286010 272856
rect 288162 272912 288218 272921
rect 288162 272847 288218 272856
rect 290922 272912 290978 272921
rect 290922 272847 290924 272856
rect 290976 272847 290978 272856
rect 293314 272912 293370 272921
rect 293314 272847 293370 272856
rect 295890 272912 295892 272921
rect 295944 272912 295946 272921
rect 295890 272847 295946 272856
rect 290924 272818 290976 272824
rect 293328 272814 293356 272847
rect 293316 272808 293368 272814
rect 293316 272750 293368 272756
rect 300858 272776 300914 272785
rect 300858 272711 300860 272720
rect 300912 272711 300914 272720
rect 303434 272776 303490 272785
rect 303434 272711 303490 272720
rect 300860 272682 300912 272688
rect 303448 272678 303476 272711
rect 303436 272672 303488 272678
rect 303436 272614 303488 272620
rect 310978 272640 311034 272649
rect 310978 272575 310980 272584
rect 311032 272575 311034 272584
rect 320914 272640 320970 272649
rect 320914 272575 320970 272584
rect 310980 272546 311032 272552
rect 320928 272542 320956 272575
rect 320916 272536 320968 272542
rect 320916 272478 320968 272484
rect 265162 272232 265218 272241
rect 265162 272167 265218 272176
rect 263598 271824 263654 271833
rect 263598 271759 263654 271768
rect 263612 271522 263640 271759
rect 263600 271516 263652 271522
rect 263600 271458 263652 271464
rect 260838 271416 260894 271425
rect 260838 271351 260840 271360
rect 260892 271351 260894 271360
rect 260840 271322 260892 271328
rect 258262 271280 258318 271289
rect 258262 271215 258318 271224
rect 264978 271280 265034 271289
rect 264978 271215 264980 271224
rect 258276 271182 258304 271215
rect 265032 271215 265034 271224
rect 264980 271186 265032 271192
rect 258264 271176 258316 271182
rect 247038 271144 247094 271153
rect 247038 271079 247094 271088
rect 252558 271144 252614 271153
rect 252558 271079 252614 271088
rect 255318 271144 255374 271153
rect 258264 271118 258316 271124
rect 255318 271079 255320 271088
rect 247052 270978 247080 271079
rect 252572 271046 252600 271079
rect 255372 271079 255374 271088
rect 255320 271050 255372 271056
rect 252560 271040 252612 271046
rect 252560 270982 252612 270988
rect 247040 270972 247092 270978
rect 247040 270914 247092 270920
rect 253938 270872 253994 270881
rect 253938 270807 253994 270816
rect 244370 270736 244426 270745
rect 244370 270671 244426 270680
rect 251270 270736 251326 270745
rect 251270 270671 251326 270680
rect 235998 270600 236054 270609
rect 235998 270535 236054 270544
rect 237378 270600 237434 270609
rect 237378 270535 237434 270544
rect 242898 270600 242954 270609
rect 242898 270535 242954 270544
rect 244278 270600 244334 270609
rect 244278 270535 244334 270544
rect 236012 268802 236040 270535
rect 237392 269754 237420 270535
rect 237380 269748 237432 269754
rect 237380 269690 237432 269696
rect 242912 268938 242940 270535
rect 244292 270298 244320 270535
rect 244280 270292 244332 270298
rect 244280 270234 244332 270240
rect 242900 268932 242952 268938
rect 242900 268874 242952 268880
rect 244384 268870 244412 270671
rect 245658 270600 245714 270609
rect 245658 270535 245714 270544
rect 247038 270600 247094 270609
rect 247038 270535 247094 270544
rect 248510 270600 248566 270609
rect 248510 270535 248566 270544
rect 249798 270600 249854 270609
rect 249798 270535 249854 270544
rect 251178 270600 251234 270609
rect 251178 270535 251234 270544
rect 245672 270434 245700 270535
rect 247052 270502 247080 270535
rect 247040 270496 247092 270502
rect 247040 270438 247092 270444
rect 245660 270428 245712 270434
rect 245660 270370 245712 270376
rect 248524 270230 248552 270535
rect 249812 270366 249840 270535
rect 249800 270360 249852 270366
rect 249800 270302 249852 270308
rect 248512 270224 248564 270230
rect 248512 270166 248564 270172
rect 251192 270162 251220 270535
rect 251180 270156 251232 270162
rect 251180 270098 251232 270104
rect 251284 269618 251312 270671
rect 252558 270600 252614 270609
rect 252558 270535 252614 270544
rect 252572 270094 252600 270535
rect 252560 270088 252612 270094
rect 252560 270030 252612 270036
rect 251272 269612 251324 269618
rect 251272 269554 251324 269560
rect 253952 269006 253980 270807
rect 255318 270736 255374 270745
rect 255318 270671 255374 270680
rect 259550 270736 259606 270745
rect 259550 270671 259606 270680
rect 253940 269000 253992 269006
rect 253940 268942 253992 268948
rect 244372 268864 244424 268870
rect 244372 268806 244424 268812
rect 236000 268796 236052 268802
rect 236000 268738 236052 268744
rect 232504 268728 232556 268734
rect 232504 268670 232556 268676
rect 230480 268660 230532 268666
rect 230480 268602 230532 268608
rect 229744 268592 229796 268598
rect 229744 268534 229796 268540
rect 220820 252544 220872 252550
rect 220820 252486 220872 252492
rect 229756 252482 229784 268534
rect 229744 252476 229796 252482
rect 229744 252418 229796 252424
rect 230492 251870 230520 268602
rect 232516 252550 232544 268670
rect 255332 268462 255360 270671
rect 256698 270600 256754 270609
rect 256698 270535 256754 270544
rect 258078 270600 258134 270609
rect 258078 270535 258134 270544
rect 259458 270600 259514 270609
rect 259458 270535 259514 270544
rect 256712 268530 256740 270535
rect 258092 269074 258120 270535
rect 258080 269068 258132 269074
rect 258080 269010 258132 269016
rect 259472 268734 259500 270535
rect 259460 268728 259512 268734
rect 259460 268670 259512 268676
rect 259564 268666 259592 270671
rect 260838 270600 260894 270609
rect 260838 270535 260894 270544
rect 262218 270600 262274 270609
rect 262218 270535 262274 270544
rect 263598 270600 263654 270609
rect 263598 270535 263654 270544
rect 259552 268660 259604 268666
rect 259552 268602 259604 268608
rect 260852 268598 260880 270535
rect 262232 269686 262260 270535
rect 263612 270026 263640 270535
rect 263600 270020 263652 270026
rect 263600 269962 263652 269968
rect 265176 269958 265204 272167
rect 276020 271924 276072 271930
rect 276020 271866 276072 271872
rect 276032 271833 276060 271866
rect 343548 271856 343600 271862
rect 270498 271824 270554 271833
rect 270498 271759 270554 271768
rect 271878 271824 271934 271833
rect 271878 271759 271934 271768
rect 276018 271824 276074 271833
rect 276018 271759 276074 271768
rect 277950 271824 278006 271833
rect 277950 271759 278006 271768
rect 280158 271824 280214 271833
rect 280158 271759 280214 271768
rect 307758 271824 307814 271833
rect 307758 271759 307760 271768
rect 270512 271726 270540 271759
rect 270500 271720 270552 271726
rect 270500 271662 270552 271668
rect 267830 271416 267886 271425
rect 267830 271351 267886 271360
rect 267844 271318 267872 271351
rect 267832 271312 267884 271318
rect 267832 271254 267884 271260
rect 266358 270600 266414 270609
rect 266358 270535 266414 270544
rect 268198 270600 268254 270609
rect 268198 270535 268254 270544
rect 265164 269952 265216 269958
rect 265164 269894 265216 269900
rect 266372 269890 266400 270535
rect 266360 269884 266412 269890
rect 266360 269826 266412 269832
rect 262220 269680 262272 269686
rect 262220 269622 262272 269628
rect 260840 268592 260892 268598
rect 260840 268534 260892 268540
rect 256700 268524 256752 268530
rect 256700 268466 256752 268472
rect 255320 268456 255372 268462
rect 255320 268398 255372 268404
rect 268212 268394 268240 270535
rect 271892 269822 271920 271759
rect 276020 271584 276072 271590
rect 276018 271552 276020 271561
rect 276072 271552 276074 271561
rect 276018 271487 276074 271496
rect 277964 271454 277992 271759
rect 280172 271658 280200 271759
rect 307812 271759 307814 271768
rect 343546 271824 343548 271833
rect 343600 271824 343602 271833
rect 343546 271759 343602 271768
rect 307760 271730 307812 271736
rect 280160 271652 280212 271658
rect 280160 271594 280212 271600
rect 277952 271448 278004 271454
rect 277952 271390 278004 271396
rect 343546 271416 343602 271425
rect 343546 271351 343602 271360
rect 343560 271318 343588 271351
rect 343548 271312 343600 271318
rect 275926 271280 275982 271289
rect 275926 271215 275982 271224
rect 278686 271280 278742 271289
rect 343548 271254 343600 271260
rect 278686 271215 278688 271224
rect 275940 271182 275968 271215
rect 278740 271215 278742 271224
rect 278688 271186 278740 271192
rect 356624 271182 356652 378150
rect 275928 271176 275980 271182
rect 356612 271176 356664 271182
rect 275928 271118 275980 271124
rect 313278 271144 313334 271153
rect 356612 271118 356664 271124
rect 313278 271079 313334 271088
rect 313292 270910 313320 271079
rect 313280 270904 313332 270910
rect 280066 270872 280122 270881
rect 313280 270846 313332 270852
rect 280066 270807 280122 270816
rect 280080 270502 280108 270807
rect 280068 270496 280120 270502
rect 280068 270438 280120 270444
rect 356612 270496 356664 270502
rect 356612 270438 356664 270444
rect 271880 269816 271932 269822
rect 271880 269758 271932 269764
rect 268200 268388 268252 268394
rect 268200 268330 268252 268336
rect 340788 253904 340840 253910
rect 340788 253846 340840 253852
rect 340800 253473 340828 253846
rect 340786 253464 340842 253473
rect 340786 253399 340842 253408
rect 339408 253292 339460 253298
rect 339408 253234 339460 253240
rect 339420 253065 339448 253234
rect 351828 253224 351880 253230
rect 351826 253192 351828 253201
rect 351880 253192 351882 253201
rect 351826 253127 351882 253136
rect 339406 253056 339462 253065
rect 339406 252991 339462 253000
rect 232504 252544 232556 252550
rect 232504 252486 232556 252492
rect 230480 251864 230532 251870
rect 230480 251806 230532 251812
rect 220820 166796 220872 166802
rect 220820 166738 220872 166744
rect 220832 145897 220860 166738
rect 260932 166728 260984 166734
rect 260932 166670 260984 166676
rect 288070 166696 288126 166705
rect 260944 166433 260972 166670
rect 265900 166660 265952 166666
rect 288070 166631 288126 166640
rect 288254 166696 288310 166705
rect 288254 166631 288310 166640
rect 291014 166696 291070 166705
rect 291014 166631 291070 166640
rect 265900 166602 265952 166608
rect 265912 166433 265940 166602
rect 285956 166456 286008 166462
rect 260930 166424 260986 166433
rect 260930 166359 260986 166368
rect 265898 166424 265954 166433
rect 288084 166433 288112 166631
rect 288268 166598 288296 166631
rect 288256 166592 288308 166598
rect 288256 166534 288308 166540
rect 291028 166530 291056 166631
rect 291016 166524 291068 166530
rect 291016 166466 291068 166472
rect 285956 166398 286008 166404
rect 288070 166424 288126 166433
rect 265898 166359 265954 166368
rect 285968 166297 285996 166398
rect 288070 166359 288126 166368
rect 293314 166424 293370 166433
rect 293314 166359 293316 166368
rect 293368 166359 293370 166368
rect 298466 166424 298522 166433
rect 298466 166359 298522 166368
rect 293316 166330 293368 166336
rect 298480 166326 298508 166359
rect 298468 166320 298520 166326
rect 285954 166288 286010 166297
rect 298468 166262 298520 166268
rect 285954 166223 286010 166232
rect 236090 165608 236146 165617
rect 236090 165543 236146 165552
rect 238758 165608 238814 165617
rect 238758 165543 238814 165552
rect 242898 165608 242954 165617
rect 242898 165543 242954 165552
rect 247130 165608 247186 165617
rect 247130 165543 247186 165552
rect 255318 165608 255374 165617
rect 255318 165543 255374 165552
rect 258170 165608 258226 165617
rect 258170 165543 258226 165552
rect 260838 165608 260894 165617
rect 260838 165543 260894 165552
rect 277398 165608 277454 165617
rect 277398 165543 277454 165552
rect 280158 165608 280214 165617
rect 280158 165543 280214 165552
rect 283378 165608 283434 165617
rect 283378 165543 283434 165552
rect 300858 165608 300914 165617
rect 300858 165543 300914 165552
rect 308218 165608 308274 165617
rect 308218 165543 308274 165552
rect 320914 165608 320970 165617
rect 320914 165543 320970 165552
rect 325882 165608 325938 165617
rect 325882 165543 325884 165552
rect 235998 164248 236054 164257
rect 235998 164183 236054 164192
rect 235264 161492 235316 161498
rect 235264 161434 235316 161440
rect 235276 146198 235304 161434
rect 236012 146266 236040 164183
rect 236104 164082 236132 165543
rect 237378 164248 237434 164257
rect 237378 164183 237434 164192
rect 236092 164076 236144 164082
rect 236092 164018 236144 164024
rect 236000 146260 236052 146266
rect 236000 146202 236052 146208
rect 235264 146192 235316 146198
rect 235264 146134 235316 146140
rect 224224 145920 224276 145926
rect 220818 145888 220874 145897
rect 224224 145862 224276 145868
rect 220818 145823 220874 145832
rect 224236 145654 224264 145862
rect 224224 145648 224276 145654
rect 224224 145590 224276 145596
rect 224316 145648 224368 145654
rect 224316 145590 224368 145596
rect 224328 145042 224356 145590
rect 236104 145518 236132 164018
rect 236644 161560 236696 161566
rect 236644 161502 236696 161508
rect 236656 146266 236684 161502
rect 236644 146260 236696 146266
rect 236644 146202 236696 146208
rect 237392 145625 237420 164183
rect 238772 148646 238800 165543
rect 240138 164248 240194 164257
rect 240138 164183 240194 164192
rect 241518 164248 241574 164257
rect 241518 164183 241574 164192
rect 238760 148640 238812 148646
rect 238760 148582 238812 148588
rect 240152 148578 240180 164183
rect 240140 148572 240192 148578
rect 240140 148514 240192 148520
rect 241532 148510 241560 164183
rect 241520 148504 241572 148510
rect 241520 148446 241572 148452
rect 242912 145722 242940 165543
rect 247038 164928 247094 164937
rect 247038 164863 247094 164872
rect 247052 164694 247080 164863
rect 247040 164688 247092 164694
rect 247040 164630 247092 164636
rect 244278 164384 244334 164393
rect 244278 164319 244334 164328
rect 244292 145926 244320 164319
rect 244370 164248 244426 164257
rect 244370 164183 244426 164192
rect 245658 164248 245714 164257
rect 245658 164183 245714 164192
rect 244280 145920 244332 145926
rect 244280 145862 244332 145868
rect 242900 145716 242952 145722
rect 242900 145658 242952 145664
rect 244384 145654 244412 164183
rect 245672 145790 245700 164183
rect 247144 145858 247172 165543
rect 255332 164966 255360 165543
rect 255320 164960 255372 164966
rect 249798 164928 249854 164937
rect 249798 164863 249800 164872
rect 249852 164863 249854 164872
rect 252558 164928 252614 164937
rect 255320 164902 255372 164908
rect 258078 164928 258134 164937
rect 252558 164863 252614 164872
rect 258078 164863 258134 164872
rect 249800 164834 249852 164840
rect 252572 164762 252600 164863
rect 258092 164830 258120 164863
rect 258080 164824 258132 164830
rect 258080 164766 258132 164772
rect 252560 164756 252612 164762
rect 252560 164698 252612 164704
rect 251270 164384 251326 164393
rect 251270 164319 251326 164328
rect 248418 164248 248474 164257
rect 248418 164183 248474 164192
rect 249890 164248 249946 164257
rect 249890 164183 249946 164192
rect 251178 164248 251234 164257
rect 251178 164183 251234 164192
rect 247132 145852 247184 145858
rect 247132 145794 247184 145800
rect 245660 145784 245712 145790
rect 245660 145726 245712 145732
rect 244372 145648 244424 145654
rect 237378 145616 237434 145625
rect 244372 145590 244424 145596
rect 248432 145586 248460 164183
rect 249904 146062 249932 164183
rect 251192 146130 251220 164183
rect 251180 146124 251232 146130
rect 251180 146066 251232 146072
rect 249892 146056 249944 146062
rect 249892 145998 249944 146004
rect 251284 145994 251312 164319
rect 252650 164248 252706 164257
rect 252650 164183 252706 164192
rect 253938 164248 253994 164257
rect 253938 164183 253994 164192
rect 255410 164248 255466 164257
rect 255410 164183 255466 164192
rect 256698 164248 256754 164257
rect 256698 164183 256754 164192
rect 251272 145988 251324 145994
rect 251272 145930 251324 145936
rect 237378 145551 237434 145560
rect 248420 145580 248472 145586
rect 248420 145522 248472 145528
rect 236092 145512 236144 145518
rect 236092 145454 236144 145460
rect 252664 145382 252692 164183
rect 253952 145450 253980 164183
rect 255424 146198 255452 164183
rect 256712 146266 256740 164183
rect 258184 162654 258212 165543
rect 259550 164384 259606 164393
rect 259550 164319 259606 164328
rect 259458 164248 259514 164257
rect 259458 164183 259514 164192
rect 259472 162790 259500 164183
rect 259460 162784 259512 162790
rect 259460 162726 259512 162732
rect 259564 162722 259592 164319
rect 260852 162858 260880 165543
rect 277412 165306 277440 165543
rect 280172 165374 280200 165543
rect 280160 165368 280212 165374
rect 280160 165310 280212 165316
rect 277400 165300 277452 165306
rect 277400 165242 277452 165248
rect 283392 165238 283420 165543
rect 300872 165442 300900 165543
rect 300860 165436 300912 165442
rect 300860 165378 300912 165384
rect 283380 165232 283432 165238
rect 264978 165200 265034 165209
rect 264978 165135 265034 165144
rect 267738 165200 267794 165209
rect 267738 165135 267740 165144
rect 263506 164248 263562 164257
rect 263782 164248 263838 164257
rect 263562 164206 263640 164234
rect 263506 164183 263562 164192
rect 260840 162852 260892 162858
rect 260840 162794 260892 162800
rect 259552 162716 259604 162722
rect 259552 162658 259604 162664
rect 258172 162648 258224 162654
rect 258172 162590 258224 162596
rect 256700 146260 256752 146266
rect 256700 146202 256752 146208
rect 255412 146192 255464 146198
rect 255412 146134 255464 146140
rect 263612 146033 263640 164206
rect 264992 164218 265020 165135
rect 267792 165135 267794 165144
rect 271878 165200 271934 165209
rect 271878 165135 271934 165144
rect 274822 165200 274878 165209
rect 274822 165135 274878 165144
rect 276018 165200 276074 165209
rect 276018 165135 276074 165144
rect 280066 165200 280122 165209
rect 283380 165174 283432 165180
rect 280066 165135 280122 165144
rect 267740 165106 267792 165112
rect 267646 164384 267702 164393
rect 267702 164342 267872 164370
rect 267646 164319 267702 164328
rect 266358 164248 266414 164257
rect 263782 164183 263838 164192
rect 264980 164212 265032 164218
rect 263796 164150 263824 164183
rect 266358 164183 266414 164192
rect 267738 164248 267794 164257
rect 267738 164183 267794 164192
rect 264980 164154 265032 164160
rect 263784 164144 263836 164150
rect 263784 164086 263836 164092
rect 266372 162178 266400 164183
rect 266360 162172 266412 162178
rect 266360 162114 266412 162120
rect 263598 146024 263654 146033
rect 263598 145959 263654 145968
rect 267752 145897 267780 164183
rect 267844 146169 267872 164342
rect 269118 164248 269174 164257
rect 269118 164183 269174 164192
rect 270498 164248 270554 164257
rect 270498 164183 270554 164192
rect 269132 146305 269160 164183
rect 270512 148442 270540 164183
rect 270500 148436 270552 148442
rect 270500 148378 270552 148384
rect 271892 148374 271920 165135
rect 273442 165064 273498 165073
rect 273442 164999 273444 165008
rect 273496 164999 273498 165008
rect 273444 164970 273496 164976
rect 273810 164384 273866 164393
rect 273810 164319 273866 164328
rect 273824 163538 273852 164319
rect 274546 164248 274602 164257
rect 274602 164206 274680 164234
rect 274546 164183 274602 164192
rect 273812 163532 273864 163538
rect 273812 163474 273864 163480
rect 274652 157334 274680 164206
rect 274652 157306 274772 157334
rect 274744 149054 274772 157306
rect 274732 149048 274784 149054
rect 274732 148990 274784 148996
rect 271880 148368 271932 148374
rect 271880 148310 271932 148316
rect 269118 146296 269174 146305
rect 274836 146266 274864 165135
rect 276032 165102 276060 165135
rect 276020 165096 276072 165102
rect 276020 165038 276072 165044
rect 277306 164248 277362 164257
rect 278042 164248 278098 164257
rect 277362 164206 277440 164234
rect 277306 164183 277362 164192
rect 277412 148986 277440 164206
rect 278042 164183 278098 164192
rect 278056 149025 278084 164183
rect 278042 149016 278098 149025
rect 277400 148980 277452 148986
rect 278042 148951 278098 148960
rect 278686 149016 278742 149025
rect 278686 148951 278742 148960
rect 277400 148922 277452 148928
rect 278700 148345 278728 148951
rect 278686 148336 278742 148345
rect 278686 148271 278742 148280
rect 269118 146231 269174 146240
rect 274824 146260 274876 146266
rect 274824 146202 274876 146208
rect 267830 146160 267886 146169
rect 267830 146095 267886 146104
rect 267738 145888 267794 145897
rect 267738 145823 267794 145832
rect 280080 145586 280108 165135
rect 308232 163985 308260 165543
rect 320928 165510 320956 165543
rect 325936 165543 325938 165552
rect 343270 165608 343326 165617
rect 343270 165543 343272 165552
rect 325884 165514 325936 165520
rect 343324 165543 343326 165552
rect 343454 165608 343510 165617
rect 343454 165543 343510 165552
rect 343272 165514 343324 165520
rect 320916 165504 320968 165510
rect 320916 165446 320968 165452
rect 343468 164898 343496 165543
rect 343456 164892 343508 164898
rect 343456 164834 343508 164840
rect 308218 163976 308274 163985
rect 308218 163911 308274 163920
rect 338488 146192 338540 146198
rect 338488 146134 338540 146140
rect 280068 145580 280120 145586
rect 280068 145522 280120 145528
rect 307668 145580 307720 145586
rect 307668 145522 307720 145528
rect 253940 145444 253992 145450
rect 253940 145386 253992 145392
rect 252652 145376 252704 145382
rect 252652 145318 252704 145324
rect 224316 145036 224368 145042
rect 224316 144978 224368 144984
rect 307680 144906 307708 145522
rect 338500 144945 338528 146134
rect 340236 146124 340288 146130
rect 340236 146066 340288 146072
rect 340248 144945 340276 146066
rect 351644 145580 351696 145586
rect 351644 145522 351696 145528
rect 351656 144945 351684 145522
rect 338486 144936 338542 144945
rect 307668 144900 307720 144906
rect 338486 144871 338542 144880
rect 340234 144936 340290 144945
rect 340234 144871 340290 144880
rect 351642 144936 351698 144945
rect 356624 144906 356652 270438
rect 356716 166734 356744 485522
rect 358268 485512 358320 485518
rect 358268 485454 358320 485460
rect 358176 485240 358228 485246
rect 358176 485182 358228 485188
rect 356888 484084 356940 484090
rect 356888 484026 356940 484032
rect 356796 468784 356848 468790
rect 356796 468726 356848 468732
rect 356808 273086 356836 468726
rect 356900 374950 356928 484026
rect 357072 475856 357124 475862
rect 357072 475798 357124 475804
rect 356980 466540 357032 466546
rect 356980 466482 357032 466488
rect 356888 374944 356940 374950
rect 356888 374886 356940 374892
rect 356992 364334 357020 466482
rect 357084 378146 357112 475798
rect 357164 473204 357216 473210
rect 357164 473146 357216 473152
rect 357072 378140 357124 378146
rect 357072 378082 357124 378088
rect 357176 376038 357204 473146
rect 358084 470484 358136 470490
rect 358084 470426 358136 470432
rect 357992 467628 358044 467634
rect 357992 467570 358044 467576
rect 357900 465588 357952 465594
rect 357900 465530 357952 465536
rect 357912 417450 357940 465530
rect 357900 417444 357952 417450
rect 357900 417386 357952 417392
rect 357532 378412 357584 378418
rect 357532 378354 357584 378360
rect 357440 378276 357492 378282
rect 357440 378218 357492 378224
rect 357164 376032 357216 376038
rect 357164 375974 357216 375980
rect 357164 375420 357216 375426
rect 357164 375362 357216 375368
rect 356992 364306 357112 364334
rect 357084 359582 357112 364306
rect 357072 359576 357124 359582
rect 357072 359518 357124 359524
rect 356796 273080 356848 273086
rect 356796 273022 356848 273028
rect 356796 271924 356848 271930
rect 356796 271866 356848 271872
rect 356808 271318 356836 271866
rect 356796 271312 356848 271318
rect 356848 271260 357020 271266
rect 356796 271254 357020 271260
rect 356808 271238 357020 271254
rect 356796 271176 356848 271182
rect 356796 271118 356848 271124
rect 356704 166728 356756 166734
rect 356704 166670 356756 166676
rect 356704 164892 356756 164898
rect 356704 164834 356756 164840
rect 351642 144871 351698 144880
rect 356612 144900 356664 144906
rect 307668 144842 307720 144848
rect 356612 144842 356664 144848
rect 235998 59800 236054 59809
rect 235998 59735 236054 59744
rect 237102 59800 237158 59809
rect 237102 59735 237158 59744
rect 255870 59800 255926 59809
rect 255870 59735 255926 59744
rect 256974 59800 257030 59809
rect 256974 59735 257030 59744
rect 262862 59800 262918 59809
rect 262862 59735 262918 59744
rect 236012 59702 236040 59735
rect 236000 59696 236052 59702
rect 236000 59638 236052 59644
rect 237116 59634 237144 59735
rect 237104 59628 237156 59634
rect 237104 59570 237156 59576
rect 255884 59566 255912 59735
rect 255872 59560 255924 59566
rect 255872 59502 255924 59508
rect 256988 59498 257016 59735
rect 260654 59664 260710 59673
rect 260654 59599 260710 59608
rect 256976 59492 257028 59498
rect 256976 59434 257028 59440
rect 259458 59392 259514 59401
rect 259458 59327 259514 59336
rect 259472 59226 259500 59327
rect 259460 59220 259512 59226
rect 259460 59162 259512 59168
rect 260668 58614 260696 59599
rect 262876 59430 262904 59735
rect 308494 59664 308550 59673
rect 308494 59599 308550 59608
rect 315854 59664 315910 59673
rect 315854 59599 315910 59608
rect 262864 59424 262916 59430
rect 261666 59392 261722 59401
rect 262864 59366 262916 59372
rect 261666 59327 261722 59336
rect 261680 59158 261708 59327
rect 279238 59256 279294 59265
rect 279238 59191 279294 59200
rect 290922 59256 290978 59265
rect 290922 59191 290978 59200
rect 300858 59256 300914 59265
rect 300858 59191 300914 59200
rect 279252 59158 279280 59191
rect 261668 59152 261720 59158
rect 261668 59094 261720 59100
rect 279240 59152 279292 59158
rect 279240 59094 279292 59100
rect 290936 59090 290964 59191
rect 290924 59084 290976 59090
rect 290924 59026 290976 59032
rect 300872 59022 300900 59191
rect 300860 59016 300912 59022
rect 300860 58958 300912 58964
rect 308508 58886 308536 59599
rect 315868 58954 315896 59599
rect 320914 59256 320970 59265
rect 320914 59191 320970 59200
rect 325882 59256 325938 59265
rect 325882 59191 325938 59200
rect 315856 58948 315908 58954
rect 315856 58890 315908 58896
rect 308496 58880 308548 58886
rect 308496 58822 308548 58828
rect 320928 58818 320956 59191
rect 320916 58812 320968 58818
rect 320916 58754 320968 58760
rect 325896 58750 325924 59191
rect 356624 59158 356652 144842
rect 356612 59152 356664 59158
rect 356612 59094 356664 59100
rect 325884 58744 325936 58750
rect 325884 58686 325936 58692
rect 260656 58608 260708 58614
rect 260656 58550 260708 58556
rect 323308 57928 323360 57934
rect 237378 57896 237434 57905
rect 237378 57831 237434 57840
rect 239218 57896 239274 57905
rect 239218 57831 239274 57840
rect 240138 57896 240194 57905
rect 240138 57831 240194 57840
rect 241610 57896 241666 57905
rect 241610 57831 241666 57840
rect 242898 57896 242954 57905
rect 242898 57831 242954 57840
rect 244370 57896 244426 57905
rect 244370 57831 244426 57840
rect 245290 57896 245346 57905
rect 245290 57831 245346 57840
rect 245658 57896 245714 57905
rect 245658 57831 245714 57840
rect 247682 57896 247738 57905
rect 247682 57831 247738 57840
rect 248418 57896 248474 57905
rect 248418 57831 248474 57840
rect 250074 57896 250130 57905
rect 250074 57831 250130 57840
rect 250994 57896 251050 57905
rect 250994 57831 251050 57840
rect 264978 57896 265034 57905
rect 264978 57831 265034 57840
rect 271050 57896 271106 57905
rect 271050 57831 271106 57840
rect 271878 57896 271934 57905
rect 271878 57831 271934 57840
rect 273258 57896 273314 57905
rect 273258 57831 273314 57840
rect 274638 57896 274694 57905
rect 274638 57831 274694 57840
rect 276938 57896 276994 57905
rect 276938 57831 276994 57840
rect 287610 57896 287666 57905
rect 287610 57831 287666 57840
rect 293314 57896 293370 57905
rect 293314 57831 293370 57840
rect 295890 57896 295946 57905
rect 295890 57831 295946 57840
rect 298098 57896 298154 57905
rect 298098 57831 298154 57840
rect 303434 57896 303490 57905
rect 303434 57831 303490 57840
rect 305826 57896 305882 57905
rect 305826 57831 305882 57840
rect 310978 57896 311034 57905
rect 310978 57831 311034 57840
rect 313370 57896 313426 57905
rect 313370 57831 313372 57840
rect 219992 56568 220044 56574
rect 219992 56510 220044 56516
rect 219900 56296 219952 56302
rect 219900 56238 219952 56244
rect 219716 54868 219768 54874
rect 219716 54810 219768 54816
rect 219256 54732 219308 54738
rect 219256 54674 219308 54680
rect 217140 54664 217192 54670
rect 217140 54606 217192 54612
rect 216496 54528 216548 54534
rect 216496 54470 216548 54476
rect 237392 54398 237420 57831
rect 239232 55894 239260 57831
rect 239220 55888 239272 55894
rect 239220 55830 239272 55836
rect 237380 54392 237432 54398
rect 237380 54334 237432 54340
rect 240152 54330 240180 57831
rect 241624 55826 241652 57831
rect 241612 55820 241664 55826
rect 241612 55762 241664 55768
rect 242912 54534 242940 57831
rect 244384 54602 244412 57831
rect 245304 55962 245332 57831
rect 245292 55956 245344 55962
rect 245292 55898 245344 55904
rect 245672 55214 245700 57831
rect 247696 56030 247724 57831
rect 247684 56024 247736 56030
rect 247684 55966 247736 55972
rect 245660 55208 245712 55214
rect 245660 55150 245712 55156
rect 248432 54670 248460 57831
rect 250088 56166 250116 57831
rect 251008 57497 251036 57831
rect 258354 57760 258410 57769
rect 258354 57695 258410 57704
rect 263598 57760 263654 57769
rect 263598 57695 263654 57704
rect 250994 57488 251050 57497
rect 250994 57423 251050 57432
rect 251178 57488 251234 57497
rect 251178 57423 251234 57432
rect 251914 57488 251970 57497
rect 251914 57423 251970 57432
rect 252558 57488 252614 57497
rect 252558 57423 252614 57432
rect 253938 57488 253994 57497
rect 253938 57423 253994 57432
rect 250076 56160 250128 56166
rect 250076 56102 250128 56108
rect 251192 54738 251220 57423
rect 251928 56098 251956 57423
rect 251916 56092 251968 56098
rect 251916 56034 251968 56040
rect 252572 54806 252600 57423
rect 253952 54874 253980 57423
rect 258368 57254 258396 57695
rect 258356 57248 258408 57254
rect 258356 57190 258408 57196
rect 263612 54942 263640 57695
rect 264992 55010 265020 57831
rect 266450 57760 266506 57769
rect 266450 57695 266506 57704
rect 268474 57760 268530 57769
rect 268474 57695 268530 57704
rect 269118 57760 269174 57769
rect 269118 57695 269174 57704
rect 266358 57488 266414 57497
rect 266358 57423 266414 57432
rect 266372 56234 266400 57423
rect 266360 56228 266412 56234
rect 266360 56170 266412 56176
rect 266464 55078 266492 57695
rect 268488 56302 268516 57695
rect 268476 56296 268528 56302
rect 268476 56238 268528 56244
rect 266452 55072 266504 55078
rect 269132 55049 269160 57695
rect 271064 56370 271092 57831
rect 271052 56364 271104 56370
rect 271052 56306 271104 56312
rect 271892 55146 271920 57831
rect 273272 56506 273300 57831
rect 273350 57760 273406 57769
rect 273350 57695 273406 57704
rect 273260 56500 273312 56506
rect 273260 56442 273312 56448
rect 271880 55140 271932 55146
rect 271880 55082 271932 55088
rect 266452 55014 266504 55020
rect 269118 55040 269174 55049
rect 264980 55004 265032 55010
rect 269118 54975 269174 54984
rect 264980 54946 265032 54952
rect 263600 54936 263652 54942
rect 263600 54878 263652 54884
rect 253940 54868 253992 54874
rect 253940 54810 253992 54816
rect 252560 54800 252612 54806
rect 252560 54742 252612 54748
rect 251180 54732 251232 54738
rect 251180 54674 251232 54680
rect 248420 54664 248472 54670
rect 248420 54606 248472 54612
rect 244372 54596 244424 54602
rect 244372 54538 244424 54544
rect 242900 54528 242952 54534
rect 242900 54470 242952 54476
rect 273364 54466 273392 57695
rect 274652 55185 274680 57831
rect 276952 56438 276980 57831
rect 287624 57322 287652 57831
rect 293328 57458 293356 57831
rect 295904 57526 295932 57831
rect 295892 57520 295944 57526
rect 295892 57462 295944 57468
rect 293316 57452 293368 57458
rect 293316 57394 293368 57400
rect 298112 57390 298140 57831
rect 303448 57662 303476 57831
rect 303436 57656 303488 57662
rect 303436 57598 303488 57604
rect 305840 57594 305868 57831
rect 310992 57730 311020 57831
rect 313424 57831 313426 57840
rect 318246 57896 318302 57905
rect 318246 57831 318302 57840
rect 323306 57896 323308 57905
rect 343180 57928 343232 57934
rect 323360 57896 323362 57905
rect 323306 57831 323362 57840
rect 343178 57896 343180 57905
rect 343232 57896 343234 57905
rect 343178 57831 343234 57840
rect 343454 57896 343510 57905
rect 356716 57866 356744 164834
rect 356808 146266 356836 271118
rect 356992 165646 357020 271238
rect 357084 253978 357112 359518
rect 357176 270502 357204 375362
rect 357452 271250 357480 378218
rect 357544 358902 357572 378354
rect 358004 374814 358032 467570
rect 358096 411942 358124 470426
rect 358084 411936 358136 411942
rect 358084 411878 358136 411884
rect 358084 390516 358136 390522
rect 358084 390458 358136 390464
rect 357992 374808 358044 374814
rect 357992 374750 358044 374756
rect 358096 359514 358124 390458
rect 358084 359508 358136 359514
rect 358084 359450 358136 359456
rect 357532 358896 357584 358902
rect 357532 358838 357584 358844
rect 358096 282198 358124 359450
rect 358084 282192 358136 282198
rect 358084 282134 358136 282140
rect 357440 271244 357492 271250
rect 357440 271186 357492 271192
rect 357164 270496 357216 270502
rect 357164 270438 357216 270444
rect 357072 253972 357124 253978
rect 357072 253914 357124 253920
rect 357256 165844 357308 165850
rect 357256 165786 357308 165792
rect 356980 165640 357032 165646
rect 356980 165582 357032 165588
rect 357268 164898 357296 165786
rect 357256 164892 357308 164898
rect 357256 164834 357308 164840
rect 357452 149025 357480 271186
rect 357624 253972 357676 253978
rect 357624 253914 357676 253920
rect 357532 165640 357584 165646
rect 357532 165582 357584 165588
rect 357438 149016 357494 149025
rect 357438 148951 357494 148960
rect 356796 146260 356848 146266
rect 356796 146202 356848 146208
rect 357544 57934 357572 165582
rect 357636 146130 357664 253914
rect 358096 253230 358124 282134
rect 358084 253224 358136 253230
rect 358084 253166 358136 253172
rect 358096 175982 358124 253166
rect 358084 175976 358136 175982
rect 358084 175918 358136 175924
rect 357624 146124 357676 146130
rect 357624 146066 357676 146072
rect 358096 145586 358124 175918
rect 358084 145580 358136 145586
rect 358084 145522 358136 145528
rect 358084 68196 358136 68202
rect 358084 68138 358136 68144
rect 358096 59362 358124 68138
rect 358084 59356 358136 59362
rect 358084 59298 358136 59304
rect 358188 58886 358216 485182
rect 358280 166802 358308 485454
rect 358360 485444 358412 485450
rect 358360 485386 358412 485392
rect 358372 166870 358400 485386
rect 363604 485376 363656 485382
rect 363604 485318 363656 485324
rect 360844 485172 360896 485178
rect 360844 485114 360896 485120
rect 359832 482860 359884 482866
rect 359832 482802 359884 482808
rect 358636 481296 358688 481302
rect 358636 481238 358688 481244
rect 358452 471368 358504 471374
rect 358452 471310 358504 471316
rect 358464 273018 358492 471310
rect 358544 468716 358596 468722
rect 358544 468658 358596 468664
rect 358452 273012 358504 273018
rect 358452 272954 358504 272960
rect 358556 271182 358584 468658
rect 358648 380526 358676 481238
rect 359464 481228 359516 481234
rect 359464 481170 359516 481176
rect 358728 477352 358780 477358
rect 358728 477294 358780 477300
rect 358636 380520 358688 380526
rect 358636 380462 358688 380468
rect 358636 378412 358688 378418
rect 358636 378354 358688 378360
rect 358648 378214 358676 378354
rect 358636 378208 358688 378214
rect 358636 378150 358688 378156
rect 358740 378078 358768 477294
rect 358820 465112 358872 465118
rect 358820 465054 358872 465060
rect 358832 460193 358860 465054
rect 358818 460184 358874 460193
rect 358818 460119 358874 460128
rect 358728 378072 358780 378078
rect 358728 378014 358780 378020
rect 358832 364334 358860 460119
rect 358910 400344 358966 400353
rect 358910 400279 358966 400288
rect 358924 369170 358952 400279
rect 359002 398168 359058 398177
rect 359002 398103 359058 398112
rect 359016 370530 359044 398103
rect 359094 394088 359150 394097
rect 359094 394023 359150 394032
rect 359004 370524 359056 370530
rect 359004 370466 359056 370472
rect 359016 369238 359044 370466
rect 359004 369232 359056 369238
rect 359004 369174 359056 369180
rect 358912 369164 358964 369170
rect 358912 369106 358964 369112
rect 358832 364306 358952 364334
rect 358636 358896 358688 358902
rect 358636 358838 358688 358844
rect 358648 271862 358676 358838
rect 358924 353161 358952 364306
rect 359108 363662 359136 394023
rect 359372 378344 359424 378350
rect 359372 378286 359424 378292
rect 359096 363656 359148 363662
rect 359096 363598 359148 363604
rect 358910 353152 358966 353161
rect 358910 353087 358966 353096
rect 358818 291816 358874 291825
rect 358818 291751 358874 291760
rect 358636 271856 358688 271862
rect 358636 271798 358688 271804
rect 358544 271176 358596 271182
rect 358544 271118 358596 271124
rect 358832 184929 358860 291751
rect 358924 246265 358952 353087
rect 359108 287609 359136 363598
rect 359188 362432 359240 362438
rect 359188 362374 359240 362380
rect 359200 362234 359228 362374
rect 359188 362228 359240 362234
rect 359188 362170 359240 362176
rect 359200 291009 359228 362170
rect 359278 292768 359334 292777
rect 359278 292703 359334 292712
rect 359186 291000 359242 291009
rect 359186 290935 359242 290944
rect 359094 287600 359150 287609
rect 359094 287535 359150 287544
rect 359108 277394 359136 287535
rect 359016 277366 359136 277394
rect 358910 246256 358966 246265
rect 358910 246191 358966 246200
rect 358818 184920 358874 184929
rect 358818 184855 358874 184864
rect 358360 166864 358412 166870
rect 358360 166806 358412 166812
rect 358268 166796 358320 166802
rect 358268 166738 358320 166744
rect 358728 145580 358780 145586
rect 358728 145522 358780 145528
rect 358740 68338 358768 145522
rect 358924 139369 358952 246191
rect 359016 180713 359044 277366
rect 359200 183433 359228 290935
rect 359292 186425 359320 292703
rect 359384 271930 359412 378286
rect 359476 377670 359504 481170
rect 359648 480140 359700 480146
rect 359648 480082 359700 480088
rect 359556 471232 359608 471238
rect 359556 471174 359608 471180
rect 359568 378826 359596 471174
rect 359660 391950 359688 480082
rect 359740 469192 359792 469198
rect 359740 469134 359792 469140
rect 359648 391944 359700 391950
rect 359648 391886 359700 391892
rect 359752 389162 359780 469134
rect 359844 414730 359872 482802
rect 360752 474360 360804 474366
rect 360752 474302 360804 474308
rect 360660 470552 360712 470558
rect 360660 470494 360712 470500
rect 359924 470416 359976 470422
rect 359924 470358 359976 470364
rect 359832 414724 359884 414730
rect 359832 414666 359884 414672
rect 359936 409154 359964 470358
rect 360016 470348 360068 470354
rect 360016 470290 360068 470296
rect 360028 410582 360056 470290
rect 360016 410576 360068 410582
rect 360016 410518 360068 410524
rect 359924 409148 359976 409154
rect 359924 409090 359976 409096
rect 359830 396808 359886 396817
rect 359830 396743 359886 396752
rect 359740 389156 359792 389162
rect 359740 389098 359792 389104
rect 359556 378820 359608 378826
rect 359556 378762 359608 378768
rect 359464 377664 359516 377670
rect 359464 377606 359516 377612
rect 359844 373994 359872 396743
rect 359922 395312 359978 395321
rect 359922 395247 359978 395256
rect 359660 373966 359872 373994
rect 359660 371890 359688 373966
rect 359936 373318 359964 395247
rect 360672 380594 360700 470494
rect 360660 380588 360712 380594
rect 360660 380530 360712 380536
rect 360764 380254 360792 474302
rect 360752 380248 360804 380254
rect 360752 380190 360804 380196
rect 359924 373312 359976 373318
rect 359924 373254 359976 373260
rect 359936 371929 359964 373254
rect 359738 371920 359794 371929
rect 359648 371884 359700 371890
rect 359738 371855 359794 371864
rect 359922 371920 359978 371929
rect 359922 371855 359978 371864
rect 359648 371826 359700 371832
rect 359464 369232 359516 369238
rect 359464 369174 359516 369180
rect 359476 291825 359504 369174
rect 359556 369164 359608 369170
rect 359556 369106 359608 369112
rect 359568 366382 359596 369106
rect 359556 366376 359608 366382
rect 359556 366318 359608 366324
rect 359568 292777 359596 366318
rect 359660 362438 359688 371826
rect 359648 362432 359700 362438
rect 359648 362374 359700 362380
rect 359554 292768 359610 292777
rect 359554 292703 359610 292712
rect 359462 291816 359518 291825
rect 359462 291751 359518 291760
rect 359752 288833 359780 371855
rect 360200 359304 360252 359310
rect 360200 359246 360252 359252
rect 360212 358834 360240 359246
rect 360200 358828 360252 358834
rect 360200 358770 360252 358776
rect 359738 288824 359794 288833
rect 359738 288759 359794 288768
rect 359752 277394 359780 288759
rect 359568 277366 359780 277394
rect 359372 271924 359424 271930
rect 359372 271866 359424 271872
rect 359278 186416 359334 186425
rect 359278 186351 359334 186360
rect 359462 186416 359518 186425
rect 359462 186351 359518 186360
rect 359370 184920 359426 184929
rect 359370 184855 359426 184864
rect 359186 183424 359242 183433
rect 359186 183359 359242 183368
rect 359094 182064 359150 182073
rect 359094 181999 359150 182008
rect 359002 180704 359058 180713
rect 359002 180639 359058 180648
rect 359016 179489 359044 180639
rect 359002 179480 359058 179489
rect 359002 179415 359058 179424
rect 358910 139360 358966 139369
rect 358910 139295 358966 139304
rect 359108 75449 359136 181999
rect 359200 76945 359228 183359
rect 359278 179480 359334 179489
rect 359278 179415 359334 179424
rect 359186 76936 359242 76945
rect 359186 76871 359242 76880
rect 359094 75440 359150 75449
rect 359094 75375 359150 75384
rect 359292 74089 359320 179415
rect 359384 78305 359412 184855
rect 359476 79937 359504 186351
rect 359568 182073 359596 277366
rect 360212 253298 360240 358770
rect 360292 271924 360344 271930
rect 360292 271866 360344 271872
rect 360200 253292 360252 253298
rect 360200 253234 360252 253240
rect 359554 182064 359610 182073
rect 359554 181999 359610 182008
rect 360212 146198 360240 253234
rect 360304 165850 360332 271866
rect 360292 165844 360344 165850
rect 360292 165786 360344 165792
rect 360200 146192 360252 146198
rect 360200 146134 360252 146140
rect 359462 79928 359518 79937
rect 359462 79863 359518 79872
rect 359370 78296 359426 78305
rect 359370 78231 359426 78240
rect 359278 74080 359334 74089
rect 359278 74015 359334 74024
rect 358728 68332 358780 68338
rect 358728 68274 358780 68280
rect 358740 68202 358768 68274
rect 358728 68196 358780 68202
rect 358728 68138 358780 68144
rect 360856 58954 360884 485114
rect 362224 483744 362276 483750
rect 362224 483686 362276 483692
rect 361304 482792 361356 482798
rect 361304 482734 361356 482740
rect 360936 474156 360988 474162
rect 360936 474098 360988 474104
rect 360948 165510 360976 474098
rect 361212 469056 361264 469062
rect 361212 468998 361264 469004
rect 361120 468988 361172 468994
rect 361120 468930 361172 468936
rect 361028 467424 361080 467430
rect 361028 467366 361080 467372
rect 361040 271454 361068 467366
rect 361132 272542 361160 468930
rect 361224 284306 361252 468998
rect 361316 376718 361344 482734
rect 361396 478644 361448 478650
rect 361396 478586 361448 478592
rect 361304 376712 361356 376718
rect 361304 376654 361356 376660
rect 361408 374882 361436 478586
rect 361488 478576 361540 478582
rect 361488 478518 361540 478524
rect 361500 378894 361528 478518
rect 361580 466608 361632 466614
rect 361580 466550 361632 466556
rect 361488 378888 361540 378894
rect 361488 378830 361540 378836
rect 361396 374876 361448 374882
rect 361396 374818 361448 374824
rect 361592 359310 361620 466550
rect 361580 359304 361632 359310
rect 361580 359246 361632 359252
rect 361212 284300 361264 284306
rect 361212 284242 361264 284248
rect 361120 272536 361172 272542
rect 361120 272478 361172 272484
rect 361028 271448 361080 271454
rect 361028 271390 361080 271396
rect 360936 165504 360988 165510
rect 360936 165446 360988 165452
rect 360844 58948 360896 58954
rect 360844 58890 360896 58896
rect 358176 58880 358228 58886
rect 358176 58822 358228 58828
rect 357532 57928 357584 57934
rect 357532 57870 357584 57876
rect 343454 57831 343456 57840
rect 313372 57802 313424 57808
rect 318260 57798 318288 57831
rect 343508 57831 343510 57840
rect 356704 57860 356756 57866
rect 343456 57802 343508 57808
rect 356704 57802 356756 57808
rect 318248 57792 318300 57798
rect 318248 57734 318300 57740
rect 310980 57724 311032 57730
rect 310980 57666 311032 57672
rect 305828 57588 305880 57594
rect 305828 57530 305880 57536
rect 362236 57526 362264 483686
rect 362684 482724 362736 482730
rect 362684 482666 362736 482672
rect 362500 482588 362552 482594
rect 362500 482530 362552 482536
rect 362408 476876 362460 476882
rect 362408 476818 362460 476824
rect 362316 475584 362368 475590
rect 362316 475526 362368 475532
rect 362328 70378 362356 475526
rect 362420 165578 362448 476818
rect 362512 271386 362540 482530
rect 362592 477216 362644 477222
rect 362592 477158 362644 477164
rect 362604 272610 362632 477158
rect 362696 376514 362724 482666
rect 362868 473068 362920 473074
rect 362868 473010 362920 473016
rect 362776 470076 362828 470082
rect 362776 470018 362828 470024
rect 362684 376508 362736 376514
rect 362684 376450 362736 376456
rect 362788 376242 362816 470018
rect 362880 380186 362908 473010
rect 363512 467492 363564 467498
rect 363512 467434 363564 467440
rect 362960 466472 363012 466478
rect 362960 466414 363012 466420
rect 362972 390522 363000 466414
rect 362960 390516 363012 390522
rect 362960 390458 363012 390464
rect 363524 380322 363552 467434
rect 363512 380316 363564 380322
rect 363512 380258 363564 380264
rect 362868 380180 362920 380186
rect 362868 380122 362920 380128
rect 362776 376236 362828 376242
rect 362776 376178 362828 376184
rect 362592 272604 362644 272610
rect 362592 272546 362644 272552
rect 362500 271380 362552 271386
rect 362500 271322 362552 271328
rect 362408 165572 362460 165578
rect 362408 165514 362460 165520
rect 362316 70372 362368 70378
rect 362316 70314 362368 70320
rect 363616 58750 363644 485318
rect 366456 485308 366508 485314
rect 366456 485250 366508 485256
rect 364064 482928 364116 482934
rect 364064 482870 364116 482876
rect 363696 481092 363748 481098
rect 363696 481034 363748 481040
rect 363708 165374 363736 481034
rect 363972 477148 364024 477154
rect 363972 477090 364024 477096
rect 363880 477012 363932 477018
rect 363880 476954 363932 476960
rect 363788 465792 363840 465798
rect 363788 465734 363840 465740
rect 363800 175234 363828 465734
rect 363892 271726 363920 476954
rect 363984 272814 364012 477090
rect 364076 375290 364104 482870
rect 364156 480004 364208 480010
rect 364156 479946 364208 479952
rect 364168 376582 364196 479946
rect 365076 478304 365128 478310
rect 365076 478246 365128 478252
rect 364248 475788 364300 475794
rect 364248 475730 364300 475736
rect 364156 376576 364208 376582
rect 364156 376518 364208 376524
rect 364260 376310 364288 475730
rect 364984 472796 365036 472802
rect 364984 472738 365036 472744
rect 364892 471776 364944 471782
rect 364892 471718 364944 471724
rect 364800 471164 364852 471170
rect 364800 471106 364852 471112
rect 364708 465656 364760 465662
rect 364708 465598 364760 465604
rect 364720 376446 364748 465598
rect 364812 379506 364840 471106
rect 364800 379500 364852 379506
rect 364800 379442 364852 379448
rect 364708 376440 364760 376446
rect 364708 376382 364760 376388
rect 364248 376304 364300 376310
rect 364248 376246 364300 376252
rect 364064 375284 364116 375290
rect 364064 375226 364116 375232
rect 364904 375086 364932 471718
rect 364892 375080 364944 375086
rect 364892 375022 364944 375028
rect 363972 272808 364024 272814
rect 363972 272750 364024 272756
rect 363880 271720 363932 271726
rect 363880 271662 363932 271668
rect 363788 175228 363840 175234
rect 363788 175170 363840 175176
rect 363696 165368 363748 165374
rect 363696 165310 363748 165316
rect 363604 58744 363656 58750
rect 363604 58686 363656 58692
rect 362224 57520 362276 57526
rect 362224 57462 362276 57468
rect 364996 57458 365024 472738
rect 365088 164898 365116 478246
rect 365536 477420 365588 477426
rect 365536 477362 365588 477368
rect 365444 477284 365496 477290
rect 365444 477226 365496 477232
rect 365352 477080 365404 477086
rect 365352 477022 365404 477028
rect 365168 468580 365220 468586
rect 365168 468522 365220 468528
rect 365180 166462 365208 468522
rect 365260 467356 365312 467362
rect 365260 467298 365312 467304
rect 365272 178022 365300 467298
rect 365364 272746 365392 477022
rect 365456 377874 365484 477226
rect 365548 380662 365576 477362
rect 366272 473136 366324 473142
rect 366272 473078 366324 473084
rect 366180 469124 366232 469130
rect 366180 469066 366232 469072
rect 365536 380656 365588 380662
rect 365536 380598 365588 380604
rect 366192 380390 366220 469066
rect 366180 380384 366232 380390
rect 366180 380326 366232 380332
rect 365626 379536 365682 379545
rect 365626 379471 365682 379480
rect 365534 379128 365590 379137
rect 365534 379063 365590 379072
rect 365444 377868 365496 377874
rect 365444 377810 365496 377816
rect 365352 272740 365404 272746
rect 365352 272682 365404 272688
rect 365548 270502 365576 379063
rect 365536 270496 365588 270502
rect 365536 270438 365588 270444
rect 365260 178016 365312 178022
rect 365260 177958 365312 177964
rect 365168 166456 365220 166462
rect 365168 166398 365220 166404
rect 365076 164892 365128 164898
rect 365076 164834 365128 164840
rect 365640 57866 365668 379471
rect 366284 376650 366312 473078
rect 366362 472696 366418 472705
rect 366362 472631 366418 472640
rect 366272 376644 366324 376650
rect 366272 376586 366324 376592
rect 365628 57860 365680 57866
rect 365628 57802 365680 57808
rect 364984 57452 365036 57458
rect 364984 57394 365036 57400
rect 298100 57384 298152 57390
rect 298100 57326 298152 57332
rect 287612 57316 287664 57322
rect 287612 57258 287664 57264
rect 276940 56432 276992 56438
rect 276940 56374 276992 56380
rect 274638 55176 274694 55185
rect 274638 55111 274694 55120
rect 273352 54460 273404 54466
rect 273352 54402 273404 54408
rect 214564 54324 214616 54330
rect 214564 54266 214616 54272
rect 240140 54324 240192 54330
rect 240140 54266 240192 54272
rect 136454 4040 136510 4049
rect 136454 3975 136510 3984
rect 132958 3496 133014 3505
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 125876 3460 125928 3466
rect 132958 3431 133014 3440
rect 125876 3402 125928 3408
rect 584 480 612 3402
rect 125888 480 125916 3402
rect 129370 3360 129426 3369
rect 129370 3295 129426 3304
rect 129384 480 129412 3295
rect 132972 480 133000 3431
rect 136468 480 136496 3975
rect 140042 3904 140098 3913
rect 140042 3839 140098 3848
rect 140056 480 140084 3839
rect 147126 3768 147182 3777
rect 147126 3703 147182 3712
rect 143538 3224 143594 3233
rect 143538 3159 143594 3168
rect 143552 480 143580 3159
rect 147140 480 147168 3703
rect 150622 3632 150678 3641
rect 150622 3567 150678 3576
rect 150636 480 150664 3567
rect 366376 3466 366404 472631
rect 366468 58818 366496 485250
rect 371884 485104 371936 485110
rect 371884 485046 371936 485052
rect 370412 483948 370464 483954
rect 370412 483890 370464 483896
rect 369216 483812 369268 483818
rect 369216 483754 369268 483760
rect 368296 480208 368348 480214
rect 368296 480150 368348 480156
rect 368020 479868 368072 479874
rect 368020 479810 368072 479816
rect 366732 479732 366784 479738
rect 366732 479674 366784 479680
rect 366548 479596 366600 479602
rect 366548 479538 366600 479544
rect 366560 165102 366588 479538
rect 366640 471300 366692 471306
rect 366640 471242 366692 471248
rect 366652 166326 366680 471242
rect 366744 273358 366772 479674
rect 367744 475516 367796 475522
rect 367744 475458 367796 475464
rect 367008 474496 367060 474502
rect 367008 474438 367060 474444
rect 366824 474292 366876 474298
rect 366824 474234 366876 474240
rect 366732 273352 366784 273358
rect 366732 273294 366784 273300
rect 366836 271318 366864 474234
rect 366916 467152 366968 467158
rect 366916 467094 366968 467100
rect 366928 282878 366956 467094
rect 367020 377466 367048 474438
rect 367560 470280 367612 470286
rect 367560 470222 367612 470228
rect 367572 380730 367600 470222
rect 367652 467560 367704 467566
rect 367652 467502 367704 467508
rect 367560 380724 367612 380730
rect 367560 380666 367612 380672
rect 367008 377460 367060 377466
rect 367008 377402 367060 377408
rect 367664 376378 367692 467502
rect 367652 376372 367704 376378
rect 367652 376314 367704 376320
rect 366916 282872 366968 282878
rect 366916 282814 366968 282820
rect 366824 271312 366876 271318
rect 366824 271254 366876 271260
rect 366640 166320 366692 166326
rect 366640 166262 366692 166268
rect 366548 165096 366600 165102
rect 366548 165038 366600 165044
rect 366456 58812 366508 58818
rect 366456 58754 366508 58760
rect 367756 57730 367784 475458
rect 367928 466200 367980 466206
rect 367928 466142 367980 466148
rect 367836 465928 367888 465934
rect 367836 465870 367888 465876
rect 367848 165034 367876 465870
rect 367940 166394 367968 466142
rect 368032 271794 368060 479810
rect 368112 476944 368164 476950
rect 368112 476886 368164 476892
rect 368020 271788 368072 271794
rect 368020 271730 368072 271736
rect 368124 271590 368152 476886
rect 368204 466404 368256 466410
rect 368204 466346 368256 466352
rect 368216 272678 368244 466346
rect 368308 375018 368336 480150
rect 368388 475720 368440 475726
rect 368388 475662 368440 475668
rect 368400 377602 368428 475662
rect 369124 475380 369176 475386
rect 369124 475322 369176 475328
rect 369032 468852 369084 468858
rect 369032 468794 369084 468800
rect 369044 385762 369072 468794
rect 369032 385756 369084 385762
rect 369032 385698 369084 385704
rect 368388 377596 368440 377602
rect 368388 377538 368440 377544
rect 368388 375420 368440 375426
rect 368388 375362 368440 375368
rect 368296 375012 368348 375018
rect 368296 374954 368348 374960
rect 368204 272672 368256 272678
rect 368204 272614 368256 272620
rect 368112 271584 368164 271590
rect 368112 271526 368164 271532
rect 368296 270496 368348 270502
rect 368296 270438 368348 270444
rect 368308 269958 368336 270438
rect 368296 269952 368348 269958
rect 368296 269894 368348 269900
rect 367928 166388 367980 166394
rect 367928 166330 367980 166336
rect 367836 165028 367888 165034
rect 367836 164970 367888 164976
rect 368308 147558 368336 269894
rect 368400 251938 368428 375362
rect 368388 251932 368440 251938
rect 368388 251874 368440 251880
rect 368296 147552 368348 147558
rect 368296 147494 368348 147500
rect 367744 57724 367796 57730
rect 367744 57666 367796 57672
rect 369136 57594 369164 475322
rect 369228 165442 369256 483754
rect 369676 482656 369728 482662
rect 369676 482598 369728 482604
rect 369492 482520 369544 482526
rect 369492 482462 369544 482468
rect 369308 479528 369360 479534
rect 369308 479470 369360 479476
rect 369216 165436 369268 165442
rect 369216 165378 369268 165384
rect 369320 164665 369348 479470
rect 369400 474088 369452 474094
rect 369400 474030 369452 474036
rect 369412 166258 369440 474030
rect 369504 271862 369532 482462
rect 369584 482452 369636 482458
rect 369584 482394 369636 482400
rect 369596 273154 369624 482394
rect 369688 380458 369716 482598
rect 370320 479936 370372 479942
rect 370320 479878 370372 479884
rect 369768 471980 369820 471986
rect 369768 471922 369820 471928
rect 369676 380452 369728 380458
rect 369676 380394 369728 380400
rect 369780 375222 369808 471922
rect 370228 471912 370280 471918
rect 370228 471854 370280 471860
rect 369860 380588 369912 380594
rect 369860 380530 369912 380536
rect 369872 379778 369900 380530
rect 369860 379772 369912 379778
rect 369860 379714 369912 379720
rect 369860 377664 369912 377670
rect 369860 377606 369912 377612
rect 369872 377534 369900 377606
rect 369860 377528 369912 377534
rect 369860 377470 369912 377476
rect 370240 375358 370268 471854
rect 370332 377942 370360 479878
rect 370320 377936 370372 377942
rect 370320 377878 370372 377884
rect 370424 376106 370452 483890
rect 370504 483676 370556 483682
rect 370504 483618 370556 483624
rect 370412 376100 370464 376106
rect 370412 376042 370464 376048
rect 370228 375352 370280 375358
rect 370228 375294 370280 375300
rect 369768 375216 369820 375222
rect 369768 375158 369820 375164
rect 370240 369854 370268 375294
rect 370240 369826 370452 369854
rect 370320 273488 370372 273494
rect 369766 273456 369822 273465
rect 370320 273430 370372 273436
rect 369766 273391 369822 273400
rect 369584 273148 369636 273154
rect 369584 273090 369636 273096
rect 369492 271856 369544 271862
rect 369492 271798 369544 271804
rect 369400 166252 369452 166258
rect 369400 166194 369452 166200
rect 369306 164656 369362 164665
rect 369306 164591 369362 164600
rect 369780 145625 369808 273391
rect 370332 145761 370360 273430
rect 370424 271998 370452 369826
rect 370412 271992 370464 271998
rect 370412 271934 370464 271940
rect 370318 145752 370374 145761
rect 370318 145687 370374 145696
rect 369766 145616 369822 145625
rect 369766 145551 369822 145560
rect 369124 57588 369176 57594
rect 369124 57530 369176 57536
rect 370516 57322 370544 483618
rect 370780 478372 370832 478378
rect 370780 478314 370832 478320
rect 370688 466132 370740 466138
rect 370688 466074 370740 466080
rect 370596 465860 370648 465866
rect 370596 465802 370648 465808
rect 370608 165306 370636 465802
rect 370700 166598 370728 466074
rect 370792 271658 370820 478314
rect 370872 472932 370924 472938
rect 370872 472874 370924 472880
rect 370884 273290 370912 472874
rect 371240 471844 371292 471850
rect 371240 471786 371292 471792
rect 371148 470144 371200 470150
rect 371148 470086 371200 470092
rect 370964 379772 371016 379778
rect 370964 379714 371016 379720
rect 370872 273284 370924 273290
rect 370872 273226 370924 273232
rect 370780 271652 370832 271658
rect 370780 271594 370832 271600
rect 370976 269822 371004 379714
rect 371160 379370 371188 470086
rect 371148 379364 371200 379370
rect 371148 379306 371200 379312
rect 371146 379264 371202 379273
rect 371146 379199 371202 379208
rect 371160 378729 371188 379199
rect 371146 378720 371202 378729
rect 371068 378678 371146 378706
rect 371068 270162 371096 378678
rect 371146 378655 371202 378664
rect 371146 376816 371202 376825
rect 371146 376751 371202 376760
rect 371056 270156 371108 270162
rect 371056 270098 371108 270104
rect 370964 269816 371016 269822
rect 370964 269758 371016 269764
rect 370688 166592 370740 166598
rect 370688 166534 370740 166540
rect 370596 165300 370648 165306
rect 370596 165242 370648 165248
rect 371068 147626 371096 270098
rect 371056 147620 371108 147626
rect 371056 147562 371108 147568
rect 371160 57662 371188 376751
rect 371252 375426 371280 471786
rect 371792 464364 371844 464370
rect 371792 464306 371844 464312
rect 371804 380594 371832 464306
rect 371792 380588 371844 380594
rect 371792 380530 371844 380536
rect 371606 378176 371662 378185
rect 371606 378111 371662 378120
rect 371240 375420 371292 375426
rect 371240 375362 371292 375368
rect 371516 375012 371568 375018
rect 371516 374954 371568 374960
rect 371528 373130 371556 374954
rect 371620 374354 371648 378111
rect 371792 375216 371844 375222
rect 371792 375158 371844 375164
rect 371804 374610 371832 375158
rect 371792 374604 371844 374610
rect 371792 374546 371844 374552
rect 371620 374326 371832 374354
rect 371528 373102 371740 373130
rect 371608 270292 371660 270298
rect 371608 270234 371660 270240
rect 371620 148986 371648 270234
rect 371712 269929 371740 373102
rect 371804 272134 371832 374326
rect 371792 272128 371844 272134
rect 371792 272070 371844 272076
rect 371698 269920 371754 269929
rect 371698 269855 371754 269864
rect 371700 267708 371752 267714
rect 371700 267650 371752 267656
rect 371712 162858 371740 267650
rect 371792 252476 371844 252482
rect 371792 252418 371844 252424
rect 371804 163538 371832 252418
rect 371792 163532 371844 163538
rect 371792 163474 371844 163480
rect 371700 162852 371752 162858
rect 371700 162794 371752 162800
rect 371608 148980 371660 148986
rect 371608 148922 371660 148928
rect 371896 59226 371924 485046
rect 376392 484016 376444 484022
rect 376392 483958 376444 483964
rect 372068 482384 372120 482390
rect 372068 482326 372120 482332
rect 371976 472660 372028 472666
rect 371976 472602 372028 472608
rect 371884 59220 371936 59226
rect 371884 59162 371936 59168
rect 371148 57656 371200 57662
rect 371148 57598 371200 57604
rect 371988 57390 372016 472602
rect 372080 165238 372108 482326
rect 372436 481364 372488 481370
rect 372436 481306 372488 481312
rect 372252 475652 372304 475658
rect 372252 475594 372304 475600
rect 372160 466064 372212 466070
rect 372160 466006 372212 466012
rect 372172 166666 372200 466006
rect 372264 271522 372292 475594
rect 372344 473000 372396 473006
rect 372344 472942 372396 472948
rect 372356 272950 372384 472942
rect 372448 379030 372476 481306
rect 374828 481024 374880 481030
rect 374828 480966 374880 480972
rect 373448 479800 373500 479806
rect 373448 479742 373500 479748
rect 373264 476808 373316 476814
rect 373264 476750 373316 476756
rect 372528 466336 372580 466342
rect 372528 466278 372580 466284
rect 372436 379024 372488 379030
rect 372436 378966 372488 378972
rect 372540 376174 372568 466278
rect 372804 385756 372856 385762
rect 372804 385698 372856 385704
rect 372816 377602 372844 385698
rect 373170 378992 373226 379001
rect 373170 378927 373226 378936
rect 373184 378729 373212 378927
rect 373170 378720 373226 378729
rect 373170 378655 373226 378664
rect 372804 377596 372856 377602
rect 372804 377538 372856 377544
rect 372528 376168 372580 376174
rect 372528 376110 372580 376116
rect 372528 375420 372580 375426
rect 372528 375362 372580 375368
rect 372540 375154 372568 375362
rect 372528 375148 372580 375154
rect 372528 375090 372580 375096
rect 372528 375012 372580 375018
rect 372528 374954 372580 374960
rect 372436 374944 372488 374950
rect 372436 374886 372488 374892
rect 372344 272944 372396 272950
rect 372344 272886 372396 272892
rect 372344 271992 372396 271998
rect 372344 271934 372396 271940
rect 372252 271516 372304 271522
rect 372252 271458 372304 271464
rect 372252 251932 372304 251938
rect 372252 251874 372304 251880
rect 372160 166660 372212 166666
rect 372160 166602 372212 166608
rect 372068 165232 372120 165238
rect 372068 165174 372120 165180
rect 372264 146169 372292 251874
rect 372356 162178 372384 271934
rect 372448 268394 372476 374886
rect 372540 374746 372568 374954
rect 372988 374808 373040 374814
rect 372988 374750 373040 374756
rect 372528 374740 372580 374746
rect 372528 374682 372580 374688
rect 372528 374604 372580 374610
rect 372528 374546 372580 374552
rect 372436 268388 372488 268394
rect 372436 268330 372488 268336
rect 372540 251190 372568 374546
rect 373000 269249 373028 374750
rect 373080 272128 373132 272134
rect 373080 272070 373132 272076
rect 372986 269240 373042 269249
rect 372986 269175 373042 269184
rect 372528 251184 372580 251190
rect 372528 251126 372580 251132
rect 372528 162852 372580 162858
rect 372528 162794 372580 162800
rect 372540 162722 372568 162794
rect 372528 162716 372580 162722
rect 372528 162658 372580 162664
rect 372344 162172 372396 162178
rect 372344 162114 372396 162120
rect 372436 148980 372488 148986
rect 372436 148922 372488 148928
rect 372250 146160 372306 146169
rect 372250 146095 372306 146104
rect 371976 57384 372028 57390
rect 371976 57326 372028 57332
rect 370504 57316 370556 57322
rect 370504 57258 370556 57264
rect 372448 54330 372476 148922
rect 372540 54466 372568 162658
rect 373092 148374 373120 272070
rect 373184 270298 373212 378655
rect 373172 270292 373224 270298
rect 373172 270234 373224 270240
rect 373276 165170 373304 476750
rect 373356 468512 373408 468518
rect 373356 468454 373408 468460
rect 373368 166530 373396 468454
rect 373460 272882 373488 479742
rect 373724 478440 373776 478446
rect 373724 478382 373776 478388
rect 373540 474224 373592 474230
rect 373540 474166 373592 474172
rect 373448 272876 373500 272882
rect 373448 272818 373500 272824
rect 373552 271017 373580 474166
rect 373632 467220 373684 467226
rect 373632 467162 373684 467168
rect 373644 271250 373672 467162
rect 373736 377806 373764 478382
rect 374460 474428 374512 474434
rect 374460 474370 374512 474376
rect 373816 471708 373868 471714
rect 373816 471650 373868 471656
rect 373724 377800 373776 377806
rect 373724 377742 373776 377748
rect 373828 375222 373856 471650
rect 373908 470212 373960 470218
rect 373908 470154 373960 470160
rect 373920 377262 373948 470154
rect 374368 468920 374420 468926
rect 374368 468862 374420 468868
rect 374274 381576 374330 381585
rect 374274 381511 374330 381520
rect 373908 377256 373960 377262
rect 373908 377198 373960 377204
rect 373816 375216 373868 375222
rect 373816 375158 373868 375164
rect 373828 369854 373856 375158
rect 373736 369826 373856 369854
rect 374288 369854 374316 381511
rect 374380 378010 374408 468862
rect 374368 378004 374420 378010
rect 374368 377946 374420 377952
rect 374472 377194 374500 474370
rect 374644 474020 374696 474026
rect 374644 473962 374696 473968
rect 374460 377188 374512 377194
rect 374460 377130 374512 377136
rect 374288 369826 374592 369854
rect 373632 271244 373684 271250
rect 373632 271186 373684 271192
rect 373538 271008 373594 271017
rect 373538 270943 373594 270952
rect 373538 269240 373594 269249
rect 373538 269175 373594 269184
rect 373356 166524 373408 166530
rect 373356 166466 373408 166472
rect 373264 165164 373316 165170
rect 373264 165106 373316 165112
rect 373552 162246 373580 269175
rect 373632 269136 373684 269142
rect 373632 269078 373684 269084
rect 373540 162240 373592 162246
rect 373540 162182 373592 162188
rect 373644 151814 373672 269078
rect 373736 252482 373764 369826
rect 373816 358080 373868 358086
rect 373816 358022 373868 358028
rect 373828 267034 373856 358022
rect 374564 277394 374592 369826
rect 374472 277366 374592 277394
rect 374472 273426 374500 277366
rect 374460 273420 374512 273426
rect 374460 273362 374512 273368
rect 374368 272332 374420 272338
rect 374368 272274 374420 272280
rect 373908 272060 373960 272066
rect 373908 272002 373960 272008
rect 373816 267028 373868 267034
rect 373816 266970 373868 266976
rect 373724 252476 373776 252482
rect 373724 252418 373776 252424
rect 373644 151786 373856 151814
rect 373828 149054 373856 151786
rect 373816 149048 373868 149054
rect 373816 148990 373868 148996
rect 373080 148368 373132 148374
rect 373080 148310 373132 148316
rect 373828 56098 373856 148990
rect 373920 144838 373948 272002
rect 374380 271289 374408 272274
rect 374366 271280 374422 271289
rect 374366 271215 374422 271224
rect 374380 163946 374408 271215
rect 374472 164150 374500 273362
rect 374552 268388 374604 268394
rect 374552 268330 374604 268336
rect 374460 164144 374512 164150
rect 374460 164086 374512 164092
rect 374368 163940 374420 163946
rect 374368 163882 374420 163888
rect 374564 161474 374592 268330
rect 374656 167006 374684 473962
rect 374736 465724 374788 465730
rect 374736 465666 374788 465672
rect 374644 167000 374696 167006
rect 374644 166942 374696 166948
rect 374748 164966 374776 465666
rect 374840 270978 374868 480966
rect 374920 479664 374972 479670
rect 374920 479606 374972 479612
rect 374932 271046 374960 479606
rect 376024 478236 376076 478242
rect 376024 478178 376076 478184
rect 375380 471640 375432 471646
rect 375380 471582 375432 471588
rect 375288 468648 375340 468654
rect 375288 468590 375340 468596
rect 375012 464432 375064 464438
rect 375012 464374 375064 464380
rect 375024 379642 375052 464374
rect 375194 381576 375250 381585
rect 375194 381511 375250 381520
rect 375208 380934 375236 381511
rect 375196 380928 375248 380934
rect 375196 380870 375248 380876
rect 375012 379636 375064 379642
rect 375012 379578 375064 379584
rect 375300 379370 375328 468590
rect 375392 379438 375420 471582
rect 375748 468444 375800 468450
rect 375748 468386 375800 468392
rect 375760 383654 375788 468386
rect 375668 383626 375788 383654
rect 375380 379432 375432 379438
rect 375380 379374 375432 379380
rect 375196 379364 375248 379370
rect 375196 379306 375248 379312
rect 375288 379364 375340 379370
rect 375288 379306 375340 379312
rect 375010 378856 375066 378865
rect 375010 378791 375066 378800
rect 374920 271040 374972 271046
rect 374920 270982 374972 270988
rect 374828 270972 374880 270978
rect 374828 270914 374880 270920
rect 374920 270020 374972 270026
rect 374920 269962 374972 269968
rect 374828 251184 374880 251190
rect 374828 251126 374880 251132
rect 374736 164960 374788 164966
rect 374736 164902 374788 164908
rect 374840 164218 374868 251126
rect 374828 164212 374880 164218
rect 374828 164154 374880 164160
rect 374840 163826 374868 164154
rect 374932 164014 374960 269962
rect 375024 269210 375052 378791
rect 375208 378758 375236 379306
rect 375196 378752 375248 378758
rect 375196 378694 375248 378700
rect 375208 378298 375236 378694
rect 375116 378270 375236 378298
rect 375116 272338 375144 378270
rect 375392 378162 375420 379374
rect 375472 378820 375524 378826
rect 375472 378762 375524 378768
rect 375484 378418 375512 378762
rect 375472 378412 375524 378418
rect 375472 378354 375524 378360
rect 375208 378134 375420 378162
rect 375104 272332 375156 272338
rect 375104 272274 375156 272280
rect 375012 269204 375064 269210
rect 375012 269146 375064 269152
rect 375208 267714 375236 378134
rect 375288 377460 375340 377466
rect 375288 377402 375340 377408
rect 375300 377330 375328 377402
rect 375288 377324 375340 377330
rect 375288 377266 375340 377272
rect 375196 267708 375248 267714
rect 375196 267650 375248 267656
rect 375300 252550 375328 377266
rect 375668 374882 375696 383626
rect 375932 377256 375984 377262
rect 375932 377198 375984 377204
rect 375840 375964 375892 375970
rect 375840 375906 375892 375912
rect 375656 374876 375708 374882
rect 375656 374818 375708 374824
rect 375748 269612 375800 269618
rect 375748 269554 375800 269560
rect 375656 269000 375708 269006
rect 375656 268942 375708 268948
rect 375288 252544 375340 252550
rect 375288 252486 375340 252492
rect 375196 252408 375248 252414
rect 375196 252350 375248 252356
rect 375208 248414 375236 252350
rect 375288 251864 375340 251870
rect 375288 251806 375340 251812
rect 375300 251190 375328 251806
rect 375288 251184 375340 251190
rect 375288 251126 375340 251132
rect 375208 248386 375328 248414
rect 375300 165646 375328 248386
rect 375288 165640 375340 165646
rect 375288 165582 375340 165588
rect 374920 164008 374972 164014
rect 374920 163950 374972 163956
rect 374840 163798 375144 163826
rect 374920 163532 374972 163538
rect 374920 163474 374972 163480
rect 374564 161446 374868 161474
rect 374840 151814 374868 161446
rect 374564 151786 374868 151814
rect 374564 145926 374592 151786
rect 374736 148504 374788 148510
rect 374736 148446 374788 148452
rect 374748 147626 374776 148446
rect 374828 148436 374880 148442
rect 374828 148378 374880 148384
rect 374736 147620 374788 147626
rect 374736 147562 374788 147568
rect 374748 146146 374776 147562
rect 374840 147558 374868 148378
rect 374828 147552 374880 147558
rect 374828 147494 374880 147500
rect 374656 146118 374776 146146
rect 374552 145920 374604 145926
rect 374552 145862 374604 145868
rect 374552 145784 374604 145790
rect 374552 145726 374604 145732
rect 373908 144832 373960 144838
rect 373908 144774 373960 144780
rect 374564 59634 374592 145726
rect 374552 59628 374604 59634
rect 374552 59570 374604 59576
rect 373816 56092 373868 56098
rect 373816 56034 373868 56040
rect 372528 54460 372580 54466
rect 372528 54402 372580 54408
rect 374656 54398 374684 146118
rect 374840 146010 374868 147494
rect 374748 145982 374868 146010
rect 374748 56030 374776 145982
rect 374828 145920 374880 145926
rect 374828 145862 374880 145868
rect 374736 56024 374788 56030
rect 374736 55966 374788 55972
rect 374840 54534 374868 145862
rect 374932 56370 374960 163474
rect 375012 162172 375064 162178
rect 375012 162114 375064 162120
rect 374920 56364 374972 56370
rect 374920 56306 374972 56312
rect 375024 55010 375052 162114
rect 375012 55004 375064 55010
rect 375012 54946 375064 54952
rect 375116 54942 375144 163798
rect 375196 148368 375248 148374
rect 375196 148310 375248 148316
rect 375208 55078 375236 148310
rect 375300 56438 375328 165582
rect 375668 145790 375696 268942
rect 375656 145784 375708 145790
rect 375656 145726 375708 145732
rect 375760 144634 375788 269554
rect 375852 269074 375880 375906
rect 375840 269068 375892 269074
rect 375840 269010 375892 269016
rect 375852 162790 375880 269010
rect 375944 269006 375972 377198
rect 375932 269000 375984 269006
rect 375932 268942 375984 268948
rect 375944 268734 375972 268942
rect 375932 268728 375984 268734
rect 375932 268670 375984 268676
rect 375932 267028 375984 267034
rect 375932 266970 375984 266976
rect 375944 162858 375972 266970
rect 376036 165345 376064 478178
rect 376116 475448 376168 475454
rect 376116 475390 376168 475396
rect 376022 165336 376078 165345
rect 376022 165271 376078 165280
rect 376128 164762 376156 475390
rect 376208 472864 376260 472870
rect 376208 472806 376260 472812
rect 376220 166938 376248 472806
rect 376300 467288 376352 467294
rect 376300 467230 376352 467236
rect 376312 271561 376340 467230
rect 376404 380905 376432 483958
rect 377312 483880 377364 483886
rect 377312 483822 377364 483828
rect 377220 481160 377272 481166
rect 377220 481102 377272 481108
rect 376576 480072 376628 480078
rect 376576 480014 376628 480020
rect 376390 380896 376446 380905
rect 376390 380831 376446 380840
rect 376484 379704 376536 379710
rect 376484 379646 376536 379652
rect 376392 378412 376444 378418
rect 376392 378354 376444 378360
rect 376298 271552 376354 271561
rect 376298 271487 376354 271496
rect 376404 269618 376432 378354
rect 376496 270337 376524 379646
rect 376588 379574 376616 480014
rect 377128 471572 377180 471578
rect 377128 471514 377180 471520
rect 376942 417888 376998 417897
rect 376942 417823 376998 417832
rect 376956 417450 376984 417823
rect 376944 417444 376996 417450
rect 376944 417386 376996 417392
rect 376956 402974 376984 417386
rect 377034 412040 377090 412049
rect 377034 411975 377090 411984
rect 377048 411942 377076 411975
rect 377036 411936 377088 411942
rect 377036 411878 377088 411884
rect 377034 410952 377090 410961
rect 377034 410887 377090 410896
rect 377048 410582 377076 410887
rect 377036 410576 377088 410582
rect 377036 410518 377088 410524
rect 376956 402946 377076 402974
rect 376944 391944 376996 391950
rect 376944 391886 376996 391892
rect 376956 390969 376984 391886
rect 376942 390960 376998 390969
rect 376942 390895 376998 390904
rect 376944 390516 376996 390522
rect 376944 390458 376996 390464
rect 376956 389337 376984 390458
rect 376942 389328 376998 389337
rect 376942 389263 376998 389272
rect 376944 389156 376996 389162
rect 376944 389098 376996 389104
rect 376956 389065 376984 389098
rect 376942 389056 376998 389065
rect 376942 388991 376998 389000
rect 376668 380656 376720 380662
rect 376668 380598 376720 380604
rect 376680 379710 376708 380598
rect 376668 379704 376720 379710
rect 376668 379646 376720 379652
rect 376576 379568 376628 379574
rect 376576 379510 376628 379516
rect 376482 270328 376538 270337
rect 376482 270263 376538 270272
rect 376392 269612 376444 269618
rect 376392 269554 376444 269560
rect 376496 258074 376524 270263
rect 376312 258046 376524 258074
rect 376208 166932 376260 166938
rect 376208 166874 376260 166880
rect 376116 164756 376168 164762
rect 376116 164698 376168 164704
rect 376116 164144 376168 164150
rect 376116 164086 376168 164092
rect 376128 163606 376156 164086
rect 376116 163600 376168 163606
rect 376116 163542 376168 163548
rect 375932 162852 375984 162858
rect 375932 162794 375984 162800
rect 375840 162784 375892 162790
rect 375840 162726 375892 162732
rect 375932 146124 375984 146130
rect 375932 146066 375984 146072
rect 375748 144628 375800 144634
rect 375748 144570 375800 144576
rect 375944 58614 375972 146066
rect 376024 144832 376076 144838
rect 376024 144774 376076 144780
rect 375932 58608 375984 58614
rect 375932 58550 375984 58556
rect 375288 56432 375340 56438
rect 375288 56374 375340 56380
rect 375196 55072 375248 55078
rect 375196 55014 375248 55020
rect 375104 54936 375156 54942
rect 375104 54878 375156 54884
rect 376036 54602 376064 144774
rect 376128 59430 376156 163542
rect 376312 162654 376340 258046
rect 376588 252414 376616 379510
rect 376666 375184 376722 375193
rect 376666 375119 376722 375128
rect 376576 252408 376628 252414
rect 376576 252350 376628 252356
rect 376576 162852 376628 162858
rect 376576 162794 376628 162800
rect 376300 162648 376352 162654
rect 376300 162590 376352 162596
rect 376208 162240 376260 162246
rect 376208 162182 376260 162188
rect 376116 59424 376168 59430
rect 376116 59366 376168 59372
rect 376220 59022 376248 162182
rect 376312 59158 376340 162590
rect 376484 162580 376536 162586
rect 376484 162522 376536 162528
rect 376392 145648 376444 145654
rect 376392 145590 376444 145596
rect 376404 144838 376432 145590
rect 376392 144832 376444 144838
rect 376392 144774 376444 144780
rect 376392 144696 376444 144702
rect 376392 144638 376444 144644
rect 376300 59152 376352 59158
rect 376300 59094 376352 59100
rect 376208 59016 376260 59022
rect 376208 58958 376260 58964
rect 376404 56234 376432 144638
rect 376496 59090 376524 162522
rect 376588 162518 376616 162794
rect 376576 162512 376628 162518
rect 376576 162454 376628 162460
rect 376484 59084 376536 59090
rect 376484 59026 376536 59032
rect 376588 56506 376616 162454
rect 376680 57934 376708 375119
rect 377048 369854 377076 402946
rect 377140 378350 377168 471514
rect 377232 380662 377260 481102
rect 377220 380656 377272 380662
rect 377220 380598 377272 380604
rect 377128 378344 377180 378350
rect 377128 378286 377180 378292
rect 377324 377330 377352 483822
rect 378784 482316 378836 482322
rect 378784 482258 378836 482264
rect 377956 471504 378008 471510
rect 377956 471446 378008 471452
rect 377496 470008 377548 470014
rect 377496 469950 377548 469956
rect 377508 422294 377536 469950
rect 377588 469940 377640 469946
rect 377588 469882 377640 469888
rect 377600 441614 377628 469882
rect 377600 441586 377812 441614
rect 377508 422266 377720 422294
rect 377692 416242 377720 422266
rect 377784 416945 377812 441586
rect 377770 416936 377826 416945
rect 377826 416894 377904 416922
rect 377770 416871 377826 416880
rect 377692 416214 377812 416242
rect 377678 414760 377734 414769
rect 377678 414695 377680 414704
rect 377732 414695 377734 414704
rect 377680 414666 377732 414672
rect 377586 412040 377642 412049
rect 377586 411975 377642 411984
rect 377496 410576 377548 410582
rect 377496 410518 377548 410524
rect 377402 409184 377458 409193
rect 377402 409119 377404 409128
rect 377456 409119 377458 409128
rect 377404 409090 377456 409096
rect 377404 379840 377456 379846
rect 377404 379782 377456 379788
rect 377312 377324 377364 377330
rect 377312 377266 377364 377272
rect 377220 374944 377272 374950
rect 377220 374886 377272 374892
rect 376956 369826 377076 369854
rect 376956 311001 376984 369826
rect 377036 358012 377088 358018
rect 377036 357954 377088 357960
rect 376942 310992 376998 311001
rect 376942 310927 376998 310936
rect 376956 287054 376984 310927
rect 376864 287026 376984 287054
rect 376760 282872 376812 282878
rect 376760 282814 376812 282820
rect 376772 282169 376800 282814
rect 376758 282160 376814 282169
rect 376758 282095 376814 282104
rect 376864 277394 376892 287026
rect 376944 284300 376996 284306
rect 376944 284242 376996 284248
rect 376956 284073 376984 284242
rect 376942 284064 376998 284073
rect 376942 283999 376998 284008
rect 376942 282296 376998 282305
rect 376942 282231 376998 282240
rect 376956 282198 376984 282231
rect 376944 282192 376996 282198
rect 376944 282134 376996 282140
rect 376864 277366 376984 277394
rect 376956 203969 376984 277366
rect 377048 270230 377076 357954
rect 377126 302152 377182 302161
rect 377126 302087 377182 302096
rect 377036 270224 377088 270230
rect 377036 270166 377088 270172
rect 377034 204232 377090 204241
rect 377034 204167 377090 204176
rect 376942 203960 376998 203969
rect 376942 203895 376998 203904
rect 377048 203017 377076 204167
rect 377034 203008 377090 203017
rect 377034 202943 377090 202952
rect 376942 201376 376998 201385
rect 376942 201311 376998 201320
rect 376956 180794 376984 201311
rect 376864 180766 376984 180794
rect 376864 171134 376892 180766
rect 376944 178016 376996 178022
rect 376944 177958 376996 177964
rect 376956 177041 376984 177958
rect 376942 177032 376998 177041
rect 376942 176967 376998 176976
rect 376944 175976 376996 175982
rect 376944 175918 376996 175924
rect 376956 175409 376984 175918
rect 376942 175400 376998 175409
rect 376942 175335 376998 175344
rect 376944 175228 376996 175234
rect 376944 175170 376996 175176
rect 376956 175137 376984 175170
rect 376942 175128 376998 175137
rect 376942 175063 376998 175072
rect 376864 171106 376984 171134
rect 376956 93809 376984 171106
rect 377048 95985 377076 202943
rect 377140 195265 377168 302087
rect 377232 270502 377260 374886
rect 377416 374678 377444 379782
rect 377404 374672 377456 374678
rect 377404 374614 377456 374620
rect 377310 310040 377366 310049
rect 377310 309975 377366 309984
rect 377220 270496 377272 270502
rect 377220 270438 377272 270444
rect 377324 204241 377352 309975
rect 377508 303929 377536 410518
rect 377600 305017 377628 411975
rect 377692 307873 377720 414666
rect 377784 413817 377812 416214
rect 377770 413808 377826 413817
rect 377770 413743 377826 413752
rect 377678 307864 377734 307873
rect 377678 307799 377734 307808
rect 377586 305008 377642 305017
rect 377586 304943 377642 304952
rect 377494 303920 377550 303929
rect 377494 303855 377550 303864
rect 377508 296714 377536 303855
rect 377508 296686 377628 296714
rect 377496 270496 377548 270502
rect 377496 270438 377548 270444
rect 377508 269142 377536 270438
rect 377496 269136 377548 269142
rect 377496 269078 377548 269084
rect 377404 252544 377456 252550
rect 377402 252512 377404 252521
rect 377456 252512 377458 252521
rect 377402 252447 377458 252456
rect 377416 252414 377444 252447
rect 377404 252408 377456 252414
rect 377404 252350 377456 252356
rect 377310 204232 377366 204241
rect 377310 204167 377366 204176
rect 377310 203960 377366 203969
rect 377310 203895 377366 203904
rect 377218 198792 377274 198801
rect 377218 198727 377274 198736
rect 377126 195256 377182 195265
rect 377126 195191 377182 195200
rect 377034 95976 377090 95985
rect 377034 95911 377090 95920
rect 376942 93800 376998 93809
rect 376942 93735 376998 93744
rect 377232 92857 377260 198727
rect 377324 96937 377352 203895
rect 377508 162858 377536 269078
rect 377600 197033 377628 296686
rect 377692 201385 377720 307799
rect 377784 306785 377812 413743
rect 377876 310049 377904 416894
rect 377968 409902 377996 471446
rect 377956 409896 378008 409902
rect 377956 409838 378008 409844
rect 378046 409184 378102 409193
rect 378046 409119 378102 409128
rect 377956 380724 378008 380730
rect 377956 380666 378008 380672
rect 377968 379846 377996 380666
rect 377956 379840 378008 379846
rect 377956 379782 378008 379788
rect 377956 375284 378008 375290
rect 377956 375226 378008 375232
rect 377968 374785 377996 375226
rect 377954 374776 378010 374785
rect 377954 374711 378010 374720
rect 377956 374672 378008 374678
rect 377956 374614 378008 374620
rect 377862 310040 377918 310049
rect 377862 309975 377918 309984
rect 377770 306776 377826 306785
rect 377770 306711 377826 306720
rect 377784 306374 377812 306711
rect 377784 306346 377904 306374
rect 377770 305008 377826 305017
rect 377770 304943 377826 304952
rect 377678 201376 377734 201385
rect 377678 201311 377734 201320
rect 377692 200841 377720 201311
rect 377678 200832 377734 200841
rect 377678 200767 377734 200776
rect 377784 200114 377812 304943
rect 377692 200086 377812 200114
rect 377692 198121 377720 200086
rect 377876 199889 377904 306346
rect 377968 270366 377996 374614
rect 378060 302161 378088 409119
rect 378140 375080 378192 375086
rect 378140 375022 378192 375028
rect 378152 374610 378180 375022
rect 378232 374876 378284 374882
rect 378232 374818 378284 374824
rect 378140 374604 378192 374610
rect 378140 374546 378192 374552
rect 378244 369854 378272 374818
rect 378152 369826 378272 369854
rect 378046 302152 378102 302161
rect 378046 302087 378102 302096
rect 378152 273494 378180 369826
rect 378692 358760 378744 358766
rect 378692 358702 378744 358708
rect 378140 273488 378192 273494
rect 378140 273430 378192 273436
rect 378600 273488 378652 273494
rect 378600 273430 378652 273436
rect 378612 273222 378640 273430
rect 378600 273216 378652 273222
rect 378600 273158 378652 273164
rect 378508 270496 378560 270502
rect 378704 270473 378732 358702
rect 378508 270438 378560 270444
rect 378690 270464 378746 270473
rect 378048 270428 378100 270434
rect 378048 270370 378100 270376
rect 377956 270360 378008 270366
rect 377956 270302 378008 270308
rect 377862 199880 377918 199889
rect 377862 199815 377918 199824
rect 377876 198801 377904 199815
rect 377862 198792 377918 198801
rect 377862 198727 377918 198736
rect 377678 198112 377734 198121
rect 377678 198047 377734 198056
rect 377586 197024 377642 197033
rect 377586 196959 377642 196968
rect 377496 162852 377548 162858
rect 377496 162794 377548 162800
rect 377588 146260 377640 146266
rect 377588 146202 377640 146208
rect 377404 146192 377456 146198
rect 377404 146134 377456 146140
rect 377416 144974 377444 146134
rect 377494 145616 377550 145625
rect 377494 145551 377550 145560
rect 377404 144968 377456 144974
rect 377404 144910 377456 144916
rect 377310 96928 377366 96937
rect 377310 96863 377366 96872
rect 377218 92848 377274 92857
rect 377218 92783 377274 92792
rect 376944 70372 376996 70378
rect 376944 70314 376996 70320
rect 376956 70009 376984 70314
rect 376942 70000 376998 70009
rect 376942 69935 376998 69944
rect 376942 68368 376998 68377
rect 376942 68303 376944 68312
rect 376996 68303 376998 68312
rect 376944 68274 376996 68280
rect 377508 59498 377536 145551
rect 377600 145314 377628 146202
rect 377588 145308 377640 145314
rect 377588 145250 377640 145256
rect 377496 59492 377548 59498
rect 377496 59434 377548 59440
rect 376668 57928 376720 57934
rect 376668 57870 376720 57876
rect 376576 56500 376628 56506
rect 376576 56442 376628 56448
rect 376392 56228 376444 56234
rect 376392 56170 376444 56176
rect 377600 54738 377628 145250
rect 377692 91089 377720 198047
rect 377862 197024 377918 197033
rect 377862 196959 377918 196968
rect 377770 195256 377826 195265
rect 377770 195191 377826 195200
rect 377678 91080 377734 91089
rect 377678 91015 377734 91024
rect 377784 88233 377812 195191
rect 377876 90001 377904 196959
rect 377968 146198 377996 270302
rect 378060 146266 378088 270370
rect 378416 252544 378468 252550
rect 378416 252486 378468 252492
rect 378428 252346 378456 252486
rect 378416 252340 378468 252346
rect 378416 252282 378468 252288
rect 378414 146296 378470 146305
rect 378048 146260 378100 146266
rect 378414 146231 378470 146240
rect 378048 146202 378100 146208
rect 377956 146192 378008 146198
rect 377956 146134 378008 146140
rect 377968 145994 377996 146134
rect 378428 146033 378456 146231
rect 378520 146130 378548 270438
rect 378690 270399 378746 270408
rect 378600 270224 378652 270230
rect 378600 270166 378652 270172
rect 378692 270224 378744 270230
rect 378692 270166 378744 270172
rect 378612 269890 378640 270166
rect 378600 269884 378652 269890
rect 378600 269826 378652 269832
rect 378612 146266 378640 269826
rect 378704 269210 378732 270166
rect 378692 269204 378744 269210
rect 378692 269146 378744 269152
rect 378796 165481 378824 482258
rect 434916 480962 434944 585239
rect 436112 522646 436140 604279
rect 436834 599584 436890 599593
rect 436834 599519 436890 599528
rect 436282 580544 436338 580553
rect 436282 580479 436338 580488
rect 436190 537024 436246 537033
rect 436190 536959 436246 536968
rect 436204 522850 436232 536959
rect 436296 527626 436324 580479
rect 436374 570344 436430 570353
rect 436374 570279 436430 570288
rect 436388 527746 436416 570279
rect 436466 565584 436522 565593
rect 436466 565519 436522 565528
rect 436376 527740 436428 527746
rect 436376 527682 436428 527688
rect 436296 527598 436416 527626
rect 436282 527504 436338 527513
rect 436282 527439 436338 527448
rect 436192 522844 436244 522850
rect 436192 522786 436244 522792
rect 436100 522640 436152 522646
rect 436100 522582 436152 522588
rect 436296 521286 436324 527439
rect 436388 522481 436416 527598
rect 436480 522918 436508 565519
rect 436558 556064 436614 556073
rect 436558 555999 436614 556008
rect 436572 522986 436600 555999
rect 436650 551304 436706 551313
rect 436650 551239 436706 551248
rect 436664 527898 436692 551239
rect 436742 541784 436798 541793
rect 436742 541719 436798 541728
rect 436756 528018 436784 541719
rect 436744 528012 436796 528018
rect 436744 527954 436796 527960
rect 436664 527870 436784 527898
rect 436652 527740 436704 527746
rect 436652 527682 436704 527688
rect 436560 522980 436612 522986
rect 436560 522922 436612 522928
rect 436468 522912 436520 522918
rect 436468 522854 436520 522860
rect 436664 522578 436692 527682
rect 436652 522572 436704 522578
rect 436652 522514 436704 522520
rect 436756 522510 436784 527870
rect 436848 522782 436876 599519
rect 457456 590345 457484 634782
rect 457720 634160 457772 634166
rect 457720 634102 457772 634108
rect 457536 634024 457588 634030
rect 457536 633966 457588 633972
rect 457548 609385 457576 633966
rect 457628 633888 457680 633894
rect 457628 633830 457680 633836
rect 457640 615505 457668 633830
rect 457732 621625 457760 634102
rect 494072 634098 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 494060 634092 494112 634098
rect 494060 634034 494112 634040
rect 471612 633752 471664 633758
rect 471612 633694 471664 633700
rect 471624 627980 471652 633694
rect 483204 633684 483256 633690
rect 483204 633626 483256 633632
rect 483216 627980 483244 633626
rect 494796 633616 494848 633622
rect 494796 633558 494848 633564
rect 494808 627980 494836 633558
rect 501236 633548 501288 633554
rect 501236 633490 501288 633496
rect 501248 627980 501276 633490
rect 512184 633480 512236 633486
rect 512184 633422 512236 633428
rect 512092 632256 512144 632262
rect 512092 632198 512144 632204
rect 512000 632188 512052 632194
rect 512000 632130 512052 632136
rect 465448 627972 465500 627978
rect 465198 627920 465448 627926
rect 465198 627914 465500 627920
rect 465198 627898 465488 627914
rect 477130 627872 477186 627881
rect 488722 627872 488778 627881
rect 477186 627830 477434 627858
rect 477130 627807 477186 627816
rect 506754 627872 506810 627881
rect 488778 627830 489026 627858
rect 488722 627807 488778 627816
rect 506810 627830 507058 627858
rect 506754 627807 506810 627816
rect 457718 621616 457774 621625
rect 457718 621551 457774 621560
rect 457626 615496 457682 615505
rect 457626 615431 457682 615440
rect 512012 612105 512040 632130
rect 512104 618905 512132 632198
rect 512196 625025 512224 633422
rect 580172 632528 580224 632534
rect 580172 632470 580224 632476
rect 580184 630873 580212 632470
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580264 627972 580316 627978
rect 580264 627914 580316 627920
rect 512182 625016 512238 625025
rect 512182 624951 512238 624960
rect 512090 618896 512146 618905
rect 512090 618831 512146 618840
rect 511998 612096 512054 612105
rect 511998 612031 512054 612040
rect 457534 609376 457590 609385
rect 457534 609311 457590 609320
rect 511998 605976 512054 605985
rect 511998 605911 512054 605920
rect 457626 602576 457682 602585
rect 457626 602511 457682 602520
rect 457534 596456 457590 596465
rect 457534 596391 457590 596400
rect 457442 590336 457498 590345
rect 457442 590271 457498 590280
rect 457442 584216 457498 584225
rect 457442 584151 457498 584160
rect 436928 528012 436980 528018
rect 436928 527954 436980 527960
rect 436836 522776 436888 522782
rect 436836 522718 436888 522724
rect 436744 522504 436796 522510
rect 436374 522472 436430 522481
rect 436744 522446 436796 522452
rect 436374 522407 436430 522416
rect 436940 521354 436968 527954
rect 457456 521422 457484 584151
rect 457444 521416 457496 521422
rect 457444 521358 457496 521364
rect 436928 521348 436980 521354
rect 436928 521290 436980 521296
rect 436284 521280 436336 521286
rect 436284 521222 436336 521228
rect 434904 480956 434956 480962
rect 434904 480898 434956 480904
rect 379244 478508 379296 478514
rect 379244 478450 379296 478456
rect 378876 478168 378928 478174
rect 378876 478110 378928 478116
rect 378782 165472 378838 165481
rect 378782 165407 378838 165416
rect 378888 164830 378916 478110
rect 378968 472728 379020 472734
rect 378968 472670 379020 472676
rect 378876 164824 378928 164830
rect 378876 164766 378928 164772
rect 378980 164694 379008 472670
rect 379060 466268 379112 466274
rect 379060 466210 379112 466216
rect 379072 271697 379100 466210
rect 379152 465996 379204 466002
rect 379152 465938 379204 465944
rect 379058 271688 379114 271697
rect 379058 271623 379114 271632
rect 379164 271114 379192 465938
rect 379256 376038 379284 478450
rect 457548 478145 457576 596391
rect 457640 518770 457668 602511
rect 459572 578054 460046 578082
rect 465092 578054 465842 578082
rect 470612 578054 471638 578082
rect 476132 578054 477434 578082
rect 483032 578054 483230 578082
rect 488552 578054 489670 578082
rect 459572 521490 459600 578054
rect 459560 521484 459612 521490
rect 459560 521426 459612 521432
rect 457628 518764 457680 518770
rect 457628 518706 457680 518712
rect 465092 517274 465120 578054
rect 470612 518838 470640 578054
rect 476132 518906 476160 578054
rect 476120 518900 476172 518906
rect 476120 518842 476172 518848
rect 470600 518832 470652 518838
rect 470600 518774 470652 518780
rect 465080 517268 465132 517274
rect 465080 517210 465132 517216
rect 483032 490521 483060 578054
rect 488552 517342 488580 578054
rect 495452 521558 495480 578068
rect 500972 578054 501262 578082
rect 506492 578054 507058 578082
rect 495440 521552 495492 521558
rect 495440 521494 495492 521500
rect 500972 520742 501000 578054
rect 500960 520736 501012 520742
rect 500960 520678 501012 520684
rect 488540 517336 488592 517342
rect 488540 517278 488592 517284
rect 506492 515409 506520 578054
rect 506478 515400 506534 515409
rect 506478 515335 506534 515344
rect 483018 490512 483074 490521
rect 483018 490447 483074 490456
rect 512012 487801 512040 605911
rect 512182 599856 512238 599865
rect 512182 599791 512238 599800
rect 512090 593736 512146 593745
rect 512090 593671 512146 593680
rect 511998 487792 512054 487801
rect 511998 487727 512054 487736
rect 512104 479505 512132 593671
rect 512196 517478 512224 599791
rect 512274 587616 512330 587625
rect 512274 587551 512330 587560
rect 512184 517472 512236 517478
rect 512184 517414 512236 517420
rect 512288 517410 512316 587551
rect 513010 580816 513066 580825
rect 513010 580751 513066 580760
rect 513024 579698 513052 580751
rect 513012 579692 513064 579698
rect 513012 579634 513064 579640
rect 560944 579692 560996 579698
rect 560944 579634 560996 579640
rect 512276 517404 512328 517410
rect 512276 517346 512328 517352
rect 560956 511970 560984 579634
rect 580276 577697 580304 627914
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 576124 518220 576176 518226
rect 576124 518162 576176 518168
rect 560944 511964 560996 511970
rect 560944 511906 560996 511912
rect 520924 495508 520976 495514
rect 520924 495450 520976 495456
rect 512090 479496 512146 479505
rect 512090 479431 512146 479440
rect 457534 478136 457590 478145
rect 457534 478071 457590 478080
rect 379336 471436 379388 471442
rect 379336 471378 379388 471384
rect 379348 378622 379376 471378
rect 379888 469872 379940 469878
rect 379888 469814 379940 469820
rect 379428 409896 379480 409902
rect 379428 409838 379480 409844
rect 379440 379522 379468 409838
rect 379900 383654 379928 469814
rect 498476 466608 498528 466614
rect 498474 466576 498476 466585
rect 517888 466608 517940 466614
rect 498528 466576 498530 466585
rect 498474 466511 498530 466520
rect 499762 466576 499818 466585
rect 499762 466511 499764 466520
rect 499816 466511 499818 466520
rect 510894 466576 510950 466585
rect 517888 466550 517940 466556
rect 510894 466511 510896 466520
rect 499764 466482 499816 466488
rect 510948 466511 510950 466520
rect 517520 466540 517572 466546
rect 510896 466482 510948 466488
rect 517520 466482 517572 466488
rect 379808 383626 379928 383654
rect 379610 382392 379666 382401
rect 379610 382327 379666 382336
rect 379440 379494 379560 379522
rect 379532 378826 379560 379494
rect 379520 378820 379572 378826
rect 379520 378762 379572 378768
rect 379336 378616 379388 378622
rect 379336 378558 379388 378564
rect 379520 378616 379572 378622
rect 379520 378558 379572 378564
rect 379428 378344 379480 378350
rect 379428 378286 379480 378292
rect 379244 376032 379296 376038
rect 379244 375974 379296 375980
rect 379336 374604 379388 374610
rect 379336 374546 379388 374552
rect 379244 358284 379296 358290
rect 379244 358226 379296 358232
rect 379152 271108 379204 271114
rect 379152 271050 379204 271056
rect 379256 270434 379284 358226
rect 379244 270428 379296 270434
rect 379244 270370 379296 270376
rect 379348 270314 379376 374546
rect 379440 273578 379468 378286
rect 379532 287054 379560 378558
rect 379624 375329 379652 382327
rect 379808 378962 379836 383626
rect 422852 380928 422904 380934
rect 422852 380870 422904 380876
rect 422864 380769 422892 380870
rect 421102 380760 421158 380769
rect 421102 380695 421158 380704
rect 422850 380760 422906 380769
rect 422850 380695 422906 380704
rect 430946 380760 431002 380769
rect 430946 380695 431002 380704
rect 433614 380760 433670 380769
rect 433614 380695 433670 380704
rect 436006 380760 436062 380769
rect 436006 380695 436062 380704
rect 438490 380760 438546 380769
rect 438490 380695 438546 380704
rect 440882 380760 440938 380769
rect 440882 380695 440938 380704
rect 443458 380760 443514 380769
rect 443458 380695 443514 380704
rect 408682 380624 408738 380633
rect 408682 380559 408738 380568
rect 413466 380624 413522 380633
rect 413466 380559 413522 380568
rect 419446 380624 419502 380633
rect 419446 380559 419502 380568
rect 408696 379846 408724 380559
rect 408684 379840 408736 379846
rect 408684 379782 408736 379788
rect 413480 379778 413508 380559
rect 413468 379772 413520 379778
rect 413468 379714 413520 379720
rect 419460 379710 419488 380559
rect 421116 380526 421144 380695
rect 430960 380662 430988 380695
rect 430948 380656 431000 380662
rect 430948 380598 431000 380604
rect 433628 380594 433656 380695
rect 434350 380624 434406 380633
rect 433616 380588 433668 380594
rect 434350 380559 434406 380568
rect 433616 380530 433668 380536
rect 421104 380520 421156 380526
rect 421104 380462 421156 380468
rect 419448 379704 419500 379710
rect 419448 379646 419500 379652
rect 381176 379636 381228 379642
rect 381176 379578 381228 379584
rect 426440 379636 426492 379642
rect 426440 379578 426492 379584
rect 380992 379024 381044 379030
rect 380992 378966 381044 378972
rect 379796 378956 379848 378962
rect 379796 378898 379848 378904
rect 379610 375320 379666 375329
rect 379610 375255 379666 375264
rect 379624 375086 379652 375255
rect 379612 375080 379664 375086
rect 379612 375022 379664 375028
rect 379532 287026 379652 287054
rect 379440 273550 379560 273578
rect 379532 273494 379560 273550
rect 379520 273488 379572 273494
rect 379426 273456 379482 273465
rect 379520 273430 379572 273436
rect 379426 273391 379482 273400
rect 379164 270286 379376 270314
rect 379164 268870 379192 270286
rect 379242 269920 379298 269929
rect 379242 269855 379298 269864
rect 379256 269385 379284 269855
rect 379242 269376 379298 269385
rect 379242 269311 379298 269320
rect 379152 268864 379204 268870
rect 379152 268806 379204 268812
rect 379060 267096 379112 267102
rect 379060 267038 379112 267044
rect 379072 265033 379100 267038
rect 379058 265024 379114 265033
rect 379058 264959 379114 264968
rect 378968 164688 379020 164694
rect 378968 164630 379020 164636
rect 379072 162790 379100 264959
rect 378968 162784 379020 162790
rect 378968 162726 379020 162732
rect 379060 162784 379112 162790
rect 379060 162726 379112 162732
rect 378980 161498 379008 162726
rect 378968 161492 379020 161498
rect 378968 161434 379020 161440
rect 378600 146260 378652 146266
rect 378600 146202 378652 146208
rect 378508 146124 378560 146130
rect 378508 146066 378560 146072
rect 378414 146024 378470 146033
rect 377956 145988 378008 145994
rect 377956 145930 378008 145936
rect 378048 145988 378100 145994
rect 378414 145959 378470 145968
rect 378048 145930 378100 145936
rect 377954 145888 378010 145897
rect 377954 145823 378010 145832
rect 377968 145625 377996 145823
rect 377954 145616 378010 145625
rect 377954 145551 378010 145560
rect 377862 89992 377918 90001
rect 377862 89927 377918 89936
rect 377770 88224 377826 88233
rect 377770 88159 377826 88168
rect 377588 54732 377640 54738
rect 377588 54674 377640 54680
rect 378060 54670 378088 145930
rect 378428 57254 378456 145959
rect 378784 145716 378836 145722
rect 378784 145658 378836 145664
rect 378692 145512 378744 145518
rect 378692 145454 378744 145460
rect 378704 59702 378732 145454
rect 378796 144634 378824 145658
rect 378876 145444 378928 145450
rect 378876 145386 378928 145392
rect 378784 144628 378836 144634
rect 378784 144570 378836 144576
rect 378692 59696 378744 59702
rect 378692 59638 378744 59644
rect 378416 57248 378468 57254
rect 378416 57190 378468 57196
rect 378796 55214 378824 144570
rect 378888 59770 378916 145386
rect 378876 59764 378928 59770
rect 378876 59706 378928 59712
rect 378980 59566 379008 161434
rect 378968 59560 379020 59566
rect 378968 59502 379020 59508
rect 378784 55208 378836 55214
rect 378784 55150 378836 55156
rect 379072 55146 379100 162726
rect 379164 145994 379192 268806
rect 379256 162586 379284 269311
rect 379244 162580 379296 162586
rect 379244 162522 379296 162528
rect 379336 146260 379388 146266
rect 379336 146202 379388 146208
rect 379244 146124 379296 146130
rect 379244 146066 379296 146072
rect 379152 145988 379204 145994
rect 379152 145930 379204 145936
rect 379256 56302 379284 146066
rect 379348 146062 379376 146202
rect 379336 146056 379388 146062
rect 379336 145998 379388 146004
rect 379244 56296 379296 56302
rect 379244 56238 379296 56244
rect 379348 56166 379376 145998
rect 379440 57798 379468 273391
rect 379532 267734 379560 273430
rect 379624 272066 379652 287026
rect 379612 272060 379664 272066
rect 379612 272002 379664 272008
rect 379624 270094 379652 272002
rect 379808 271153 379836 378898
rect 380900 378888 380952 378894
rect 380900 378830 380952 378836
rect 379980 378820 380032 378826
rect 379980 378762 380032 378768
rect 379888 377528 379940 377534
rect 379888 377470 379940 377476
rect 379900 377194 379928 377470
rect 379888 377188 379940 377194
rect 379888 377130 379940 377136
rect 379794 271144 379850 271153
rect 379794 271079 379850 271088
rect 379702 270464 379758 270473
rect 379702 270399 379758 270408
rect 379612 270088 379664 270094
rect 379612 270030 379664 270036
rect 379716 269793 379744 270399
rect 379808 270026 379836 271079
rect 379796 270020 379848 270026
rect 379796 269962 379848 269968
rect 379702 269784 379758 269793
rect 379702 269719 379758 269728
rect 379532 267706 379652 267734
rect 379624 171134 379652 267706
rect 379532 171106 379652 171134
rect 379532 164082 379560 171106
rect 379716 164150 379744 269719
rect 379900 269006 379928 377130
rect 379992 270502 380020 378762
rect 380912 378486 380940 378830
rect 381004 378554 381032 378966
rect 380992 378548 381044 378554
rect 380992 378490 381044 378496
rect 380900 378480 380952 378486
rect 380900 378422 380952 378428
rect 380912 377074 380940 378422
rect 381004 377210 381032 378490
rect 381004 377182 381124 377210
rect 380912 377046 381032 377074
rect 380900 376984 380952 376990
rect 380900 376926 380952 376932
rect 380912 358766 380940 376926
rect 380900 358760 380952 358766
rect 380900 358702 380952 358708
rect 381004 358018 381032 377046
rect 381096 358290 381124 377182
rect 381188 376990 381216 379578
rect 426452 379409 426480 379578
rect 434364 379574 434392 380559
rect 436020 380458 436048 380695
rect 436008 380452 436060 380458
rect 436008 380394 436060 380400
rect 438504 380390 438532 380695
rect 438492 380384 438544 380390
rect 438492 380326 438544 380332
rect 440896 380322 440924 380695
rect 440884 380316 440936 380322
rect 440884 380258 440936 380264
rect 443472 380254 443500 380695
rect 445942 380624 445998 380633
rect 445942 380559 445998 380568
rect 443460 380248 443512 380254
rect 443460 380190 443512 380196
rect 445956 380186 445984 380559
rect 445944 380180 445996 380186
rect 445944 380122 445996 380128
rect 434352 379568 434404 379574
rect 434352 379510 434404 379516
rect 439044 379500 439096 379506
rect 439044 379442 439096 379448
rect 435732 379432 435784 379438
rect 396078 379400 396134 379409
rect 396078 379335 396134 379344
rect 397090 379400 397146 379409
rect 397090 379335 397146 379344
rect 403622 379400 403678 379409
rect 403622 379335 403678 379344
rect 405830 379400 405886 379409
rect 405830 379335 405886 379344
rect 407578 379400 407634 379409
rect 407578 379335 407634 379344
rect 408314 379400 408370 379409
rect 408314 379335 408316 379344
rect 396092 378690 396120 379335
rect 397104 378962 397132 379335
rect 402978 379264 403034 379273
rect 402978 379199 403034 379208
rect 397092 378956 397144 378962
rect 397092 378898 397144 378904
rect 396080 378684 396132 378690
rect 396080 378626 396132 378632
rect 402992 377330 403020 379199
rect 403636 378826 403664 379335
rect 405370 379264 405426 379273
rect 405370 379199 405426 379208
rect 403624 378820 403676 378826
rect 403624 378762 403676 378768
rect 402980 377324 403032 377330
rect 402980 377266 403032 377272
rect 381176 376984 381228 376990
rect 381176 376926 381228 376932
rect 381176 376032 381228 376038
rect 381176 375974 381228 375980
rect 381084 358284 381136 358290
rect 381084 358226 381136 358232
rect 381188 358086 381216 375974
rect 405384 375018 405412 379199
rect 405844 378622 405872 379335
rect 405832 378616 405884 378622
rect 405832 378558 405884 378564
rect 407592 378418 407620 379335
rect 408368 379335 408370 379344
rect 411258 379400 411314 379409
rect 411258 379335 411314 379344
rect 412362 379400 412418 379409
rect 412362 379335 412418 379344
rect 413098 379400 413154 379409
rect 413098 379335 413154 379344
rect 414570 379400 414626 379409
rect 414570 379335 414626 379344
rect 423402 379400 423458 379409
rect 423402 379335 423458 379344
rect 426438 379400 426494 379409
rect 426438 379335 426494 379344
rect 426622 379400 426678 379409
rect 426622 379335 426678 379344
rect 435730 379400 435732 379409
rect 439056 379409 439084 379442
rect 435784 379400 435786 379409
rect 435730 379335 435786 379344
rect 439042 379400 439098 379409
rect 439042 379335 439098 379344
rect 447506 379400 447562 379409
rect 447506 379335 447562 379344
rect 451002 379400 451058 379409
rect 451002 379335 451058 379344
rect 452750 379400 452806 379409
rect 452750 379335 452806 379344
rect 455602 379400 455658 379409
rect 455602 379335 455658 379344
rect 458362 379400 458418 379409
rect 458362 379335 458418 379344
rect 460938 379400 460994 379409
rect 460938 379335 460994 379344
rect 463514 379400 463570 379409
rect 463514 379335 463570 379344
rect 474830 379400 474886 379409
rect 474830 379335 474886 379344
rect 408316 379306 408368 379312
rect 410062 379264 410118 379273
rect 410062 379199 410118 379208
rect 407580 378412 407632 378418
rect 407580 378354 407632 378360
rect 409970 378176 410026 378185
rect 409970 378111 410026 378120
rect 405372 375012 405424 375018
rect 405372 374954 405424 374960
rect 409984 374610 410012 378111
rect 410076 377398 410104 379199
rect 411272 378486 411300 379335
rect 412376 378554 412404 379335
rect 412364 378548 412416 378554
rect 412364 378490 412416 378496
rect 411260 378480 411312 378486
rect 411260 378422 411312 378428
rect 413112 377602 413140 379335
rect 413100 377596 413152 377602
rect 413100 377538 413152 377544
rect 414584 377534 414612 379335
rect 415766 379264 415822 379273
rect 415766 379199 415822 379208
rect 416042 379264 416098 379273
rect 416042 379199 416098 379208
rect 414572 377528 414624 377534
rect 414572 377470 414624 377476
rect 415780 377466 415808 379199
rect 415768 377460 415820 377466
rect 415768 377402 415820 377408
rect 410064 377392 410116 377398
rect 410064 377334 410116 377340
rect 416056 376106 416084 379199
rect 418250 378720 418306 378729
rect 418250 378655 418306 378664
rect 416962 378584 417018 378593
rect 416962 378519 417018 378528
rect 416044 376100 416096 376106
rect 416044 376042 416096 376048
rect 416976 375970 417004 378519
rect 418158 378176 418214 378185
rect 418158 378111 418214 378120
rect 416964 375964 417016 375970
rect 416964 375906 417016 375912
rect 418172 374950 418200 378111
rect 418264 376174 418292 378655
rect 419630 378176 419686 378185
rect 419630 378111 419686 378120
rect 421746 378176 421802 378185
rect 421746 378111 421802 378120
rect 418252 376168 418304 376174
rect 418252 376110 418304 376116
rect 418160 374944 418212 374950
rect 418160 374886 418212 374892
rect 419644 374746 419672 378111
rect 421760 374814 421788 378111
rect 423416 377670 423444 379335
rect 425978 378720 426034 378729
rect 425978 378655 426034 378664
rect 423954 378176 424010 378185
rect 423954 378111 424010 378120
rect 425150 378176 425206 378185
rect 425150 378111 425206 378120
rect 423404 377664 423456 377670
rect 423404 377606 423456 377612
rect 423968 375086 423996 378111
rect 423956 375080 424008 375086
rect 423956 375022 424008 375028
rect 425164 374882 425192 378111
rect 425992 376242 426020 378655
rect 426636 378350 426664 379335
rect 437754 379264 437810 379273
rect 437754 379199 437810 379208
rect 427910 378720 427966 378729
rect 427910 378655 427966 378664
rect 426624 378344 426676 378350
rect 426624 378286 426676 378292
rect 427924 376310 427952 378655
rect 436466 378584 436522 378593
rect 436466 378519 436522 378528
rect 431130 378312 431186 378321
rect 431130 378247 431186 378256
rect 428278 378176 428334 378185
rect 428278 378111 428334 378120
rect 429290 378176 429346 378185
rect 429290 378111 429346 378120
rect 427912 376304 427964 376310
rect 427912 376246 427964 376252
rect 425980 376236 426032 376242
rect 425980 376178 426032 376184
rect 428292 375154 428320 378111
rect 428280 375148 428332 375154
rect 428280 375090 428332 375096
rect 425152 374876 425204 374882
rect 425152 374818 425204 374824
rect 421748 374808 421800 374814
rect 421748 374750 421800 374756
rect 419632 374740 419684 374746
rect 419632 374682 419684 374688
rect 429304 374678 429332 378111
rect 431144 375358 431172 378247
rect 432234 378176 432290 378185
rect 432234 378111 432290 378120
rect 431132 375352 431184 375358
rect 431132 375294 431184 375300
rect 432248 375222 432276 378111
rect 436480 376038 436508 378519
rect 436468 376032 436520 376038
rect 436468 375974 436520 375980
rect 437768 375290 437796 379199
rect 439056 378350 439084 379335
rect 439044 378344 439096 378350
rect 439044 378286 439096 378292
rect 447520 377874 447548 379335
rect 447508 377868 447560 377874
rect 447508 377810 447560 377816
rect 451016 377738 451044 379335
rect 452764 377942 452792 379335
rect 452752 377936 452804 377942
rect 452752 377878 452804 377884
rect 455616 377806 455644 379335
rect 458376 378010 458404 379335
rect 460952 378078 460980 379335
rect 460940 378072 460992 378078
rect 463528 378049 463556 379335
rect 473450 379264 473506 379273
rect 473450 379199 473506 379208
rect 465078 379128 465134 379137
rect 465078 379063 465134 379072
rect 460940 378014 460992 378020
rect 463514 378040 463570 378049
rect 458364 378004 458416 378010
rect 463514 377975 463570 377984
rect 458364 377946 458416 377952
rect 455604 377800 455656 377806
rect 455604 377742 455656 377748
rect 451004 377732 451056 377738
rect 451004 377674 451056 377680
rect 465092 376378 465120 379063
rect 467930 378856 467986 378865
rect 467930 378791 467986 378800
rect 470874 378856 470930 378865
rect 470874 378791 470930 378800
rect 467944 376446 467972 378791
rect 470888 376514 470916 378791
rect 473464 376582 473492 379199
rect 474844 378146 474872 379335
rect 480534 379264 480590 379273
rect 480534 379199 480590 379208
rect 503074 379264 503130 379273
rect 503074 379199 503130 379208
rect 503534 379264 503590 379273
rect 503534 379199 503590 379208
rect 477590 378992 477646 379001
rect 477590 378927 477646 378936
rect 474832 378140 474884 378146
rect 474832 378082 474884 378088
rect 477604 376718 477632 378927
rect 477592 376712 477644 376718
rect 477592 376654 477644 376660
rect 480548 376650 480576 379199
rect 483386 378992 483442 379001
rect 483386 378927 483442 378936
rect 483400 376689 483428 378927
rect 503088 378282 503116 379199
rect 503076 378276 503128 378282
rect 503076 378218 503128 378224
rect 503548 378214 503576 379199
rect 516600 378344 516652 378350
rect 516600 378286 516652 378292
rect 503536 378208 503588 378214
rect 503536 378150 503588 378156
rect 483386 376680 483442 376689
rect 480536 376644 480588 376650
rect 483386 376615 483442 376624
rect 480536 376586 480588 376592
rect 473452 376576 473504 376582
rect 473452 376518 473504 376524
rect 470876 376508 470928 376514
rect 470876 376450 470928 376456
rect 467932 376440 467984 376446
rect 467932 376382 467984 376388
rect 465080 376372 465132 376378
rect 465080 376314 465132 376320
rect 437756 375284 437808 375290
rect 437756 375226 437808 375232
rect 432236 375216 432288 375222
rect 432236 375158 432288 375164
rect 429292 374672 429344 374678
rect 429292 374614 429344 374620
rect 409972 374604 410024 374610
rect 409972 374546 410024 374552
rect 500776 359712 500828 359718
rect 500776 359654 500828 359660
rect 498936 359576 498988 359582
rect 498936 359518 498988 359524
rect 498948 358873 498976 359518
rect 500788 358873 500816 359654
rect 498934 358864 498990 358873
rect 498934 358799 498990 358808
rect 500774 358864 500830 358873
rect 500774 358799 500830 358808
rect 510894 358864 510950 358873
rect 510894 358799 510896 358808
rect 510948 358799 510950 358808
rect 510896 358770 510948 358776
rect 381176 358080 381228 358086
rect 381176 358022 381228 358028
rect 380992 358012 381044 358018
rect 380992 357954 381044 357960
rect 421102 273592 421158 273601
rect 421102 273527 421158 273536
rect 422850 273592 422906 273601
rect 422850 273527 422906 273536
rect 427634 273592 427690 273601
rect 427634 273527 427690 273536
rect 445942 273592 445998 273601
rect 445942 273527 445998 273536
rect 421116 273358 421144 273527
rect 422864 273426 422892 273527
rect 427648 273494 427676 273527
rect 427636 273488 427688 273494
rect 427636 273430 427688 273436
rect 422852 273420 422904 273426
rect 422852 273362 422904 273368
rect 421104 273352 421156 273358
rect 421104 273294 421156 273300
rect 445956 273290 445984 273527
rect 445944 273284 445996 273290
rect 445944 273226 445996 273232
rect 425244 273216 425296 273222
rect 425244 273158 425296 273164
rect 423404 273148 423456 273154
rect 423404 273090 423456 273096
rect 423416 273057 423444 273090
rect 425256 273057 425284 273158
rect 425980 273080 426032 273086
rect 423402 273048 423458 273057
rect 423402 272983 423458 272992
rect 425242 273048 425298 273057
rect 425242 272983 425298 272992
rect 425978 273048 425980 273057
rect 426032 273048 426034 273057
rect 425978 272983 426034 272992
rect 428186 273048 428242 273057
rect 428186 272983 428188 272992
rect 428240 272983 428242 272992
rect 468482 273048 468538 273057
rect 468482 272983 468538 272992
rect 428188 272954 428240 272960
rect 468496 272950 468524 272983
rect 468484 272944 468536 272950
rect 468484 272886 468536 272892
rect 470874 272912 470930 272921
rect 470874 272847 470930 272856
rect 478418 272912 478474 272921
rect 478418 272847 478420 272856
rect 470888 272814 470916 272847
rect 478472 272847 478474 272856
rect 478420 272818 478472 272824
rect 470876 272808 470928 272814
rect 470876 272750 470928 272756
rect 473450 272776 473506 272785
rect 473450 272711 473452 272720
rect 473504 272711 473506 272720
rect 480810 272776 480866 272785
rect 480810 272711 480866 272720
rect 473452 272682 473504 272688
rect 480824 272678 480852 272711
rect 480812 272672 480864 272678
rect 475842 272640 475898 272649
rect 480812 272614 480864 272620
rect 485962 272640 486018 272649
rect 475842 272575 475844 272584
rect 475896 272575 475898 272584
rect 485962 272575 486018 272584
rect 475844 272546 475896 272552
rect 485976 272542 486004 272575
rect 485964 272536 486016 272542
rect 485964 272478 486016 272484
rect 401690 272232 401746 272241
rect 401690 272167 401746 272176
rect 415858 272232 415914 272241
rect 415858 272167 415914 272176
rect 416042 272232 416098 272241
rect 416042 272167 416098 272176
rect 455786 272232 455842 272241
rect 455786 272167 455842 272176
rect 396724 272060 396776 272066
rect 396724 272002 396776 272008
rect 379980 270496 380032 270502
rect 379980 270438 380032 270444
rect 379992 270026 380020 270438
rect 380440 270428 380492 270434
rect 380440 270370 380492 270376
rect 379980 270020 380032 270026
rect 379980 269962 380032 269968
rect 379980 269816 380032 269822
rect 379980 269758 380032 269764
rect 379888 269000 379940 269006
rect 379888 268942 379940 268948
rect 379704 164144 379756 164150
rect 379704 164086 379756 164092
rect 379520 164076 379572 164082
rect 379520 164018 379572 164024
rect 379428 57792 379480 57798
rect 379428 57734 379480 57740
rect 379336 56160 379388 56166
rect 379336 56102 379388 56108
rect 379060 55140 379112 55146
rect 379060 55082 379112 55088
rect 379532 54806 379560 164018
rect 379612 162852 379664 162858
rect 379612 162794 379664 162800
rect 379624 162314 379652 162794
rect 379612 162308 379664 162314
rect 379612 162250 379664 162256
rect 379624 59294 379652 162250
rect 379716 161474 379744 164086
rect 379796 162852 379848 162858
rect 379796 162794 379848 162800
rect 379808 162518 379836 162794
rect 379796 162512 379848 162518
rect 379796 162454 379848 162460
rect 379716 161446 379836 161474
rect 379612 59288 379664 59294
rect 379612 59230 379664 59236
rect 379808 54874 379836 161446
rect 379900 145382 379928 268942
rect 379992 146130 380020 269758
rect 380452 269618 380480 270370
rect 380440 269612 380492 269618
rect 380440 269554 380492 269560
rect 390558 269376 390614 269385
rect 390558 269311 390614 269320
rect 388442 269240 388498 269249
rect 388442 269175 388498 269184
rect 388456 268938 388484 269175
rect 388444 268932 388496 268938
rect 388444 268874 388496 268880
rect 390572 268802 390600 269311
rect 391940 269136 391992 269142
rect 391940 269078 391992 269084
rect 390560 268796 390612 268802
rect 390560 268738 390612 268744
rect 391952 268666 391980 269078
rect 391940 268660 391992 268666
rect 391940 268602 391992 268608
rect 396736 252414 396764 272002
rect 397458 270600 397514 270609
rect 397458 270535 397514 270544
rect 398838 270600 398894 270609
rect 398838 270535 398894 270544
rect 400218 270600 400274 270609
rect 400218 270535 400274 270544
rect 397472 270162 397500 270535
rect 397460 270156 397512 270162
rect 397460 270098 397512 270104
rect 398852 269958 398880 270535
rect 400232 270298 400260 270535
rect 400220 270292 400272 270298
rect 400220 270234 400272 270240
rect 401704 270230 401732 272167
rect 415872 272066 415900 272167
rect 415860 272060 415912 272066
rect 415860 272002 415912 272008
rect 416056 271182 416084 272167
rect 433340 272128 433392 272134
rect 433340 272070 433392 272076
rect 430580 271992 430632 271998
rect 430580 271934 430632 271940
rect 425704 271924 425756 271930
rect 425704 271866 425756 271872
rect 427820 271924 427872 271930
rect 427820 271866 427872 271872
rect 416044 271176 416096 271182
rect 409878 271144 409934 271153
rect 409878 271079 409934 271088
rect 412730 271144 412786 271153
rect 416044 271118 416096 271124
rect 418158 271144 418214 271153
rect 412730 271079 412786 271088
rect 418158 271079 418160 271088
rect 409892 270978 409920 271079
rect 412744 271046 412772 271079
rect 418212 271079 418214 271088
rect 418160 271050 418212 271056
rect 412732 271040 412784 271046
rect 412732 270982 412784 270988
rect 409880 270972 409932 270978
rect 409880 270914 409932 270920
rect 405738 270872 405794 270881
rect 405738 270807 405794 270816
rect 402978 270600 403034 270609
rect 402978 270535 403034 270544
rect 403622 270600 403678 270609
rect 403622 270535 403678 270544
rect 404358 270600 404414 270609
rect 404358 270535 404414 270544
rect 401692 270224 401744 270230
rect 401692 270166 401744 270172
rect 398840 269952 398892 269958
rect 398840 269894 398892 269900
rect 402992 268734 403020 270535
rect 403636 270026 403664 270535
rect 403624 270020 403676 270026
rect 403624 269962 403676 269968
rect 402980 268728 403032 268734
rect 402980 268670 403032 268676
rect 404372 268394 404400 270535
rect 405752 270094 405780 270807
rect 411350 270736 411406 270745
rect 411350 270671 411406 270680
rect 407118 270600 407174 270609
rect 407118 270535 407174 270544
rect 408498 270600 408554 270609
rect 408498 270535 408554 270544
rect 409878 270600 409934 270609
rect 409878 270535 409934 270544
rect 411258 270600 411314 270609
rect 411258 270535 411314 270544
rect 407132 270434 407160 270535
rect 407120 270428 407172 270434
rect 407120 270370 407172 270376
rect 408512 270366 408540 270535
rect 408500 270360 408552 270366
rect 408500 270302 408552 270308
rect 405740 270088 405792 270094
rect 405740 270030 405792 270036
rect 409892 268870 409920 270535
rect 411272 270502 411300 270535
rect 411260 270496 411312 270502
rect 411260 270438 411312 270444
rect 411364 269890 411392 270671
rect 413006 270600 413062 270609
rect 413006 270535 413062 270544
rect 414018 270600 414074 270609
rect 414018 270535 414074 270544
rect 416778 270600 416834 270609
rect 416778 270535 416834 270544
rect 418158 270600 418214 270609
rect 418158 270535 418214 270544
rect 419538 270600 419594 270609
rect 419538 270535 419594 270544
rect 420918 270600 420974 270609
rect 420918 270535 420974 270544
rect 411352 269884 411404 269890
rect 411352 269826 411404 269832
rect 413020 269822 413048 270535
rect 413008 269816 413060 269822
rect 413008 269758 413060 269764
rect 414032 269006 414060 270535
rect 416792 269074 416820 270535
rect 416780 269068 416832 269074
rect 416780 269010 416832 269016
rect 414020 269000 414072 269006
rect 414020 268942 414072 268948
rect 409880 268864 409932 268870
rect 409880 268806 409932 268812
rect 418172 268666 418200 270535
rect 419552 268802 419580 270535
rect 420932 268938 420960 270535
rect 420920 268932 420972 268938
rect 420920 268874 420972 268880
rect 419540 268796 419592 268802
rect 419540 268738 419592 268744
rect 418160 268660 418212 268666
rect 418160 268602 418212 268608
rect 404360 268388 404412 268394
rect 404360 268330 404412 268336
rect 396724 252408 396776 252414
rect 396724 252350 396776 252356
rect 425716 251938 425744 271866
rect 427832 271833 427860 271866
rect 430592 271833 430620 271934
rect 433352 271833 433380 272070
rect 427818 271824 427874 271833
rect 427818 271759 427874 271768
rect 430578 271824 430634 271833
rect 430578 271759 430634 271768
rect 432050 271824 432106 271833
rect 432050 271759 432106 271768
rect 433338 271824 433394 271833
rect 433338 271759 433394 271768
rect 434718 271824 434774 271833
rect 434718 271759 434774 271768
rect 437478 271824 437534 271833
rect 437478 271759 437534 271768
rect 442998 271824 443054 271833
rect 442998 271759 443054 271768
rect 447138 271824 447194 271833
rect 447138 271759 447194 271768
rect 449898 271824 449954 271833
rect 449898 271759 449954 271768
rect 452658 271824 452714 271833
rect 455800 271794 455828 272167
rect 458180 271856 458232 271862
rect 458178 271824 458180 271833
rect 458232 271824 458234 271833
rect 452658 271759 452714 271768
rect 455788 271788 455840 271794
rect 432064 271454 432092 271759
rect 426992 271448 427044 271454
rect 426992 271390 427044 271396
rect 427084 271448 427136 271454
rect 427084 271390 427136 271396
rect 432052 271448 432104 271454
rect 432052 271390 432104 271396
rect 433338 271416 433394 271425
rect 427004 271182 427032 271390
rect 426992 271176 427044 271182
rect 426992 271118 427044 271124
rect 427096 252482 427124 271390
rect 434732 271386 434760 271759
rect 433338 271351 433394 271360
rect 434720 271380 434772 271386
rect 433352 271182 433380 271351
rect 434720 271322 434772 271328
rect 437492 271318 437520 271759
rect 443012 271590 443040 271759
rect 443000 271584 443052 271590
rect 443000 271526 443052 271532
rect 447152 271522 447180 271759
rect 449912 271726 449940 271759
rect 449900 271720 449952 271726
rect 449900 271662 449952 271668
rect 452672 271658 452700 271759
rect 458178 271759 458234 271768
rect 455788 271730 455840 271736
rect 503626 271688 503682 271697
rect 452660 271652 452712 271658
rect 503626 271623 503682 271632
rect 452660 271594 452712 271600
rect 447140 271516 447192 271522
rect 447140 271458 447192 271464
rect 440238 271416 440294 271425
rect 503640 271386 503668 271623
rect 440238 271351 440294 271360
rect 503628 271380 503680 271386
rect 437480 271312 437532 271318
rect 437480 271254 437532 271260
rect 440146 271280 440202 271289
rect 440252 271250 440280 271351
rect 503628 271322 503680 271328
rect 503626 271280 503682 271289
rect 440146 271215 440202 271224
rect 440240 271244 440292 271250
rect 440160 271182 440188 271215
rect 503626 271215 503628 271224
rect 440240 271186 440292 271192
rect 503680 271215 503682 271224
rect 503628 271186 503680 271192
rect 516612 271182 516640 378286
rect 517532 358834 517560 466482
rect 517796 466472 517848 466478
rect 517796 466414 517848 466420
rect 517612 378276 517664 378282
rect 517612 378218 517664 378224
rect 517520 358828 517572 358834
rect 517520 358770 517572 358776
rect 433340 271176 433392 271182
rect 433340 271118 433392 271124
rect 440148 271176 440200 271182
rect 440148 271118 440200 271124
rect 516600 271176 516652 271182
rect 516600 271118 516652 271124
rect 434718 270872 434774 270881
rect 434718 270807 434774 270816
rect 436098 270872 436154 270881
rect 436098 270807 436154 270816
rect 437478 270872 437534 270881
rect 437478 270807 437534 270816
rect 429198 270736 429254 270745
rect 429198 270671 429254 270680
rect 427084 252476 427136 252482
rect 427084 252418 427136 252424
rect 425704 251932 425756 251938
rect 425704 251874 425756 251880
rect 429212 251870 429240 270671
rect 434732 252550 434760 270807
rect 434810 270736 434866 270745
rect 434810 270671 434866 270680
rect 434824 267714 434852 270671
rect 434812 267708 434864 267714
rect 434812 267650 434864 267656
rect 436112 267034 436140 270807
rect 437492 267102 437520 270807
rect 437480 267096 437532 267102
rect 437480 267038 437532 267044
rect 436100 267028 436152 267034
rect 436100 266970 436152 266976
rect 500868 253360 500920 253366
rect 500866 253328 500868 253337
rect 500920 253328 500922 253337
rect 499212 253292 499264 253298
rect 500866 253263 500922 253272
rect 499212 253234 499264 253240
rect 499224 252793 499252 253234
rect 499210 252784 499266 252793
rect 499210 252719 499266 252728
rect 510894 252648 510950 252657
rect 510894 252583 510896 252592
rect 510948 252583 510950 252592
rect 510896 252554 510948 252560
rect 434720 252544 434772 252550
rect 434720 252486 434772 252492
rect 429200 251864 429252 251870
rect 429200 251806 429252 251812
rect 428280 167000 428332 167006
rect 428280 166942 428332 166948
rect 418436 166864 418488 166870
rect 418434 166832 418436 166841
rect 428292 166841 428320 166942
rect 430948 166932 431000 166938
rect 430948 166874 431000 166880
rect 430960 166841 430988 166874
rect 418488 166832 418490 166841
rect 418434 166767 418490 166776
rect 421010 166832 421066 166841
rect 421010 166767 421012 166776
rect 421064 166767 421066 166776
rect 428278 166832 428334 166841
rect 428278 166767 428334 166776
rect 430946 166832 431002 166841
rect 430946 166767 431002 166776
rect 433614 166832 433670 166841
rect 433614 166767 433670 166776
rect 473450 166832 473506 166841
rect 473450 166767 473506 166776
rect 475842 166832 475898 166841
rect 475842 166767 475898 166776
rect 478418 166832 478474 166841
rect 478418 166767 478474 166776
rect 480902 166832 480958 166841
rect 480902 166767 480958 166776
rect 421012 166738 421064 166744
rect 433628 166734 433656 166767
rect 433616 166728 433668 166734
rect 433616 166670 433668 166676
rect 473464 166598 473492 166767
rect 475856 166666 475884 166767
rect 475844 166660 475896 166666
rect 475844 166602 475896 166608
rect 473452 166592 473504 166598
rect 434350 166560 434406 166569
rect 473452 166534 473504 166540
rect 434350 166495 434406 166504
rect 423402 166288 423458 166297
rect 423402 166223 423404 166232
rect 423456 166223 423458 166232
rect 423404 166194 423456 166200
rect 434364 165646 434392 166495
rect 478432 166462 478460 166767
rect 480916 166530 480944 166767
rect 483386 166696 483442 166705
rect 483386 166631 483442 166640
rect 485962 166696 486018 166705
rect 485962 166631 486018 166640
rect 480904 166524 480956 166530
rect 480904 166466 480956 166472
rect 478420 166456 478472 166462
rect 478420 166398 478472 166404
rect 483400 166394 483428 166631
rect 483388 166388 483440 166394
rect 483388 166330 483440 166336
rect 485976 166326 486004 166631
rect 503258 166560 503314 166569
rect 503258 166495 503314 166504
rect 485964 166320 486016 166326
rect 485964 166262 486016 166268
rect 434352 165640 434404 165646
rect 397458 165608 397514 165617
rect 397458 165543 397514 165552
rect 401598 165608 401654 165617
rect 401598 165543 401654 165552
rect 404358 165608 404414 165617
rect 404358 165543 404414 165552
rect 407118 165608 407174 165617
rect 407118 165543 407174 165552
rect 415490 165608 415546 165617
rect 415490 165543 415546 165552
rect 416042 165608 416098 165617
rect 416042 165543 416098 165552
rect 418710 165608 418766 165617
rect 418710 165543 418766 165552
rect 423678 165608 423734 165617
rect 423678 165543 423734 165552
rect 426530 165608 426586 165617
rect 426530 165543 426586 165552
rect 429658 165608 429714 165617
rect 434352 165582 434404 165588
rect 435086 165608 435142 165617
rect 429658 165543 429714 165552
rect 435086 165543 435142 165552
rect 435914 165608 435970 165617
rect 435914 165543 435970 165552
rect 437938 165608 437994 165617
rect 437938 165543 437994 165552
rect 438490 165608 438546 165617
rect 438490 165543 438546 165552
rect 440146 165608 440202 165617
rect 440146 165543 440202 165552
rect 440882 165608 440938 165617
rect 440882 165543 440938 165552
rect 443458 165608 443514 165617
rect 443458 165543 443514 165552
rect 445850 165608 445906 165617
rect 445850 165543 445906 165552
rect 447322 165608 447378 165617
rect 447322 165543 447378 165552
rect 449898 165608 449954 165617
rect 449898 165543 449954 165552
rect 452658 165608 452714 165617
rect 452658 165543 452714 165552
rect 455418 165608 455474 165617
rect 455418 165543 455474 165552
rect 458362 165608 458418 165617
rect 458362 165543 458364 165552
rect 396170 164384 396226 164393
rect 396170 164319 396226 164328
rect 396078 164248 396134 164257
rect 396078 164183 396134 164192
rect 396092 163946 396120 164183
rect 396184 164014 396212 164319
rect 396172 164008 396224 164014
rect 396172 163950 396224 163956
rect 396080 163940 396132 163946
rect 396080 163882 396132 163888
rect 379980 146124 380032 146130
rect 379980 146066 380032 146072
rect 396092 145518 396120 163882
rect 396080 145512 396132 145518
rect 396080 145454 396132 145460
rect 396184 145450 396212 163950
rect 396724 161492 396776 161498
rect 396724 161434 396776 161440
rect 396736 146198 396764 161434
rect 397472 148510 397500 165543
rect 398838 164248 398894 164257
rect 398838 164183 398894 164192
rect 400218 164248 400274 164257
rect 400218 164183 400274 164192
rect 397460 148504 397512 148510
rect 397460 148446 397512 148452
rect 398852 148442 398880 164183
rect 400232 148986 400260 164183
rect 401612 149054 401640 165543
rect 403070 164384 403126 164393
rect 403070 164319 403126 164328
rect 402978 164248 403034 164257
rect 402978 164183 403034 164192
rect 401600 149048 401652 149054
rect 401600 148990 401652 148996
rect 400220 148980 400272 148986
rect 400220 148922 400272 148928
rect 398840 148436 398892 148442
rect 398840 148378 398892 148384
rect 396724 146192 396776 146198
rect 396724 146134 396776 146140
rect 402992 145790 403020 164183
rect 403084 146266 403112 164319
rect 403072 146260 403124 146266
rect 403072 146202 403124 146208
rect 404372 145858 404400 165543
rect 407132 164694 407160 165543
rect 412638 164928 412694 164937
rect 412638 164863 412640 164872
rect 412692 164863 412694 164872
rect 412640 164834 412692 164840
rect 409878 164792 409934 164801
rect 409878 164727 409880 164736
rect 409932 164727 409934 164736
rect 409880 164698 409932 164704
rect 407120 164688 407172 164694
rect 407120 164630 407172 164636
rect 411350 164384 411406 164393
rect 411350 164319 411406 164328
rect 405738 164248 405794 164257
rect 405738 164183 405794 164192
rect 407210 164248 407266 164257
rect 407210 164183 407266 164192
rect 408498 164248 408554 164257
rect 408498 164183 408554 164192
rect 409970 164248 410026 164257
rect 409970 164183 410026 164192
rect 411258 164248 411314 164257
rect 411258 164183 411314 164192
rect 404360 145852 404412 145858
rect 404360 145794 404412 145800
rect 402980 145784 403032 145790
rect 402980 145726 403032 145732
rect 405752 145654 405780 164183
rect 407224 145722 407252 164183
rect 408512 145926 408540 164183
rect 409984 145994 410012 164183
rect 411272 146062 411300 164183
rect 411260 146056 411312 146062
rect 411260 145998 411312 146004
rect 409972 145988 410024 145994
rect 409972 145930 410024 145936
rect 408500 145920 408552 145926
rect 408500 145862 408552 145868
rect 407212 145716 407264 145722
rect 407212 145658 407264 145664
rect 405740 145648 405792 145654
rect 405740 145590 405792 145596
rect 396172 145444 396224 145450
rect 396172 145386 396224 145392
rect 379888 145376 379940 145382
rect 379888 145318 379940 145324
rect 379900 59362 379928 145318
rect 411364 145314 411392 164319
rect 412638 164248 412694 164257
rect 412638 164183 412694 164192
rect 414018 164248 414074 164257
rect 414018 164183 414074 164192
rect 412652 146130 412680 164183
rect 412640 146124 412692 146130
rect 412640 146066 412692 146072
rect 414032 145382 414060 164183
rect 415504 146033 415532 165543
rect 416056 164830 416084 165543
rect 416044 164824 416096 164830
rect 416044 164766 416096 164772
rect 416778 164248 416834 164257
rect 416778 164183 416834 164192
rect 418158 164248 418214 164257
rect 418158 164183 418214 164192
rect 416792 146198 416820 164183
rect 418172 162314 418200 164183
rect 418724 162654 418752 165543
rect 420918 164520 420974 164529
rect 420918 164455 420974 164464
rect 419538 164248 419594 164257
rect 419538 164183 419594 164192
rect 418712 162648 418764 162654
rect 418712 162590 418764 162596
rect 419552 162586 419580 164183
rect 419540 162580 419592 162586
rect 419540 162522 419592 162528
rect 418160 162308 418212 162314
rect 418160 162250 418212 162256
rect 420932 162246 420960 164455
rect 422298 164248 422354 164257
rect 422298 164183 422354 164192
rect 422312 163606 422340 164183
rect 422300 163600 422352 163606
rect 422300 163542 422352 163548
rect 420920 162240 420972 162246
rect 420920 162182 420972 162188
rect 416780 146192 416832 146198
rect 416780 146134 416832 146140
rect 415490 146024 415546 146033
rect 415490 145959 415546 145968
rect 423692 145897 423720 165543
rect 425058 164248 425114 164257
rect 425058 164183 425114 164192
rect 426438 164248 426494 164257
rect 426438 164183 426494 164192
rect 423678 145888 423734 145897
rect 423678 145823 423734 145832
rect 425072 145761 425100 164183
rect 426452 164150 426480 164183
rect 426440 164144 426492 164150
rect 426440 164086 426492 164092
rect 426544 164082 426572 165543
rect 427820 164348 427872 164354
rect 427820 164290 427872 164296
rect 426532 164076 426584 164082
rect 426532 164018 426584 164024
rect 427832 162722 427860 164290
rect 429106 164248 429162 164257
rect 429162 164206 429240 164234
rect 429672 164218 429700 165543
rect 432234 165064 432290 165073
rect 432234 164999 432290 165008
rect 430578 164520 430634 164529
rect 430578 164455 430634 164464
rect 429106 164183 429162 164192
rect 427820 162716 427872 162722
rect 427820 162658 427872 162664
rect 425058 145752 425114 145761
rect 425058 145687 425114 145696
rect 429212 145625 429240 164206
rect 429660 164212 429712 164218
rect 429660 164154 429712 164160
rect 430592 162178 430620 164455
rect 432248 163538 432276 164999
rect 435100 164354 435128 165543
rect 435928 165034 435956 165543
rect 435916 165028 435968 165034
rect 435916 164970 435968 164976
rect 436190 164928 436246 164937
rect 436190 164863 436246 164872
rect 435088 164348 435140 164354
rect 435088 164290 435140 164296
rect 434626 164248 434682 164257
rect 434682 164206 434760 164234
rect 434626 164183 434682 164192
rect 432236 163532 432288 163538
rect 432236 163474 432288 163480
rect 430580 162172 430632 162178
rect 430580 162114 430632 162120
rect 434732 148374 434760 164206
rect 436204 162858 436232 164863
rect 436192 162852 436244 162858
rect 436192 162794 436244 162800
rect 437952 162790 437980 165543
rect 438504 165102 438532 165543
rect 440160 165102 440188 165543
rect 438492 165096 438544 165102
rect 438492 165038 438544 165044
rect 440148 165096 440200 165102
rect 440148 165038 440200 165044
rect 440160 164506 440188 165038
rect 440896 164966 440924 165543
rect 443472 165374 443500 165543
rect 443460 165368 443512 165374
rect 443460 165310 443512 165316
rect 445864 165170 445892 165543
rect 447336 165238 447364 165543
rect 449912 165306 449940 165543
rect 452672 165510 452700 165543
rect 452660 165504 452712 165510
rect 452660 165446 452712 165452
rect 455432 165442 455460 165543
rect 458416 165543 458418 165552
rect 458364 165514 458416 165520
rect 455420 165436 455472 165442
rect 455420 165378 455472 165384
rect 449900 165300 449952 165306
rect 449900 165242 449952 165248
rect 447324 165232 447376 165238
rect 447324 165174 447376 165180
rect 503272 165170 503300 166495
rect 503350 165608 503406 165617
rect 503350 165543 503406 165552
rect 445852 165164 445904 165170
rect 445852 165106 445904 165112
rect 503260 165164 503312 165170
rect 503260 165106 503312 165112
rect 503364 165034 503392 165543
rect 516612 165102 516640 271118
rect 517532 252618 517560 358770
rect 517624 271386 517652 378218
rect 517704 378208 517756 378214
rect 517704 378150 517756 378156
rect 517716 271862 517744 378150
rect 517808 359650 517836 466414
rect 517796 359644 517848 359650
rect 517796 359586 517848 359592
rect 517900 359582 517928 466550
rect 518900 465112 518952 465118
rect 518900 465054 518952 465060
rect 518912 459649 518940 465054
rect 518898 459640 518954 459649
rect 518898 459575 518954 459584
rect 519450 459640 519506 459649
rect 519450 459575 519506 459584
rect 519082 400344 519138 400353
rect 519082 400279 519138 400288
rect 518990 398168 519046 398177
rect 518990 398103 519046 398112
rect 519004 369238 519032 398103
rect 518992 369232 519044 369238
rect 518992 369174 519044 369180
rect 517980 359644 518032 359650
rect 517980 359586 518032 359592
rect 517888 359576 517940 359582
rect 517888 359518 517940 359524
rect 517900 354674 517928 359518
rect 517808 354646 517928 354674
rect 517704 271856 517756 271862
rect 517704 271798 517756 271804
rect 517612 271380 517664 271386
rect 517612 271322 517664 271328
rect 517520 252612 517572 252618
rect 517520 252554 517572 252560
rect 516600 165096 516652 165102
rect 516600 165038 516652 165044
rect 503352 165028 503404 165034
rect 503352 164970 503404 164976
rect 517532 164966 517560 252554
rect 517624 165170 517652 271322
rect 517704 253360 517756 253366
rect 517704 253302 517756 253308
rect 517716 253230 517744 253302
rect 517808 253298 517836 354646
rect 517888 271856 517940 271862
rect 517888 271798 517940 271804
rect 517900 271250 517928 271798
rect 517888 271244 517940 271250
rect 517888 271186 517940 271192
rect 517796 253292 517848 253298
rect 517796 253234 517848 253240
rect 517704 253224 517756 253230
rect 517704 253166 517756 253172
rect 517612 165164 517664 165170
rect 517612 165106 517664 165112
rect 440884 164960 440936 164966
rect 440884 164902 440936 164908
rect 510528 164960 510580 164966
rect 510528 164902 510580 164908
rect 517520 164960 517572 164966
rect 517520 164902 517572 164908
rect 440160 164478 440280 164506
rect 437940 162784 437992 162790
rect 437940 162726 437992 162732
rect 434720 148368 434772 148374
rect 440252 148345 440280 164478
rect 434720 148310 434772 148316
rect 440238 148336 440294 148345
rect 440238 148271 440294 148280
rect 500224 146192 500276 146198
rect 500224 146134 500276 146140
rect 498660 146124 498712 146130
rect 498660 146066 498712 146072
rect 429198 145616 429254 145625
rect 429198 145551 429254 145560
rect 414020 145376 414072 145382
rect 414020 145318 414072 145324
rect 411352 145308 411404 145314
rect 411352 145250 411404 145256
rect 498672 144945 498700 146066
rect 500236 144945 500264 146134
rect 510540 145586 510568 164902
rect 517520 146192 517572 146198
rect 517520 146134 517572 146140
rect 517532 145654 517560 146134
rect 517520 145648 517572 145654
rect 517520 145590 517572 145596
rect 510528 145580 510580 145586
rect 510528 145522 510580 145528
rect 510540 145466 510568 145522
rect 510618 145480 510674 145489
rect 510540 145438 510618 145466
rect 510618 145415 510674 145424
rect 498658 144936 498714 144945
rect 498658 144871 498714 144880
rect 500222 144936 500278 144945
rect 500222 144871 500278 144880
rect 396078 59800 396134 59809
rect 396078 59735 396134 59744
rect 397090 59800 397146 59809
rect 397090 59735 397092 59744
rect 396092 59702 396120 59735
rect 397144 59735 397146 59744
rect 403070 59800 403126 59809
rect 403070 59735 403126 59744
rect 416962 59800 417018 59809
rect 416962 59735 417018 59744
rect 422850 59800 422906 59809
rect 422850 59735 422906 59744
rect 423954 59800 424010 59809
rect 423954 59735 424010 59744
rect 397092 59706 397144 59712
rect 396080 59696 396132 59702
rect 396080 59638 396132 59644
rect 403084 59634 403112 59735
rect 404174 59664 404230 59673
rect 403072 59628 403124 59634
rect 404174 59599 404230 59608
rect 412546 59664 412602 59673
rect 412546 59599 412602 59608
rect 403072 59570 403124 59576
rect 379888 59356 379940 59362
rect 379888 59298 379940 59304
rect 404188 58614 404216 59599
rect 410706 59392 410762 59401
rect 410706 59327 410762 59336
rect 410720 59226 410748 59327
rect 410708 59220 410760 59226
rect 410708 59162 410760 59168
rect 404176 58608 404228 58614
rect 404176 58550 404228 58556
rect 397458 57896 397514 57905
rect 397458 57831 397514 57840
rect 399482 57896 399538 57905
rect 399482 57831 399538 57840
rect 400218 57896 400274 57905
rect 400218 57831 400274 57840
rect 401690 57896 401746 57905
rect 401690 57831 401746 57840
rect 404358 57896 404414 57905
rect 404358 57831 404414 57840
rect 405830 57896 405886 57905
rect 405830 57831 405886 57840
rect 407210 57896 407266 57905
rect 407210 57831 407266 57840
rect 408314 57896 408370 57905
rect 408314 57831 408370 57840
rect 408682 57896 408738 57905
rect 408682 57831 408738 57840
rect 409878 57896 409934 57905
rect 409878 57831 409934 57840
rect 411350 57896 411406 57905
rect 411350 57831 411406 57840
rect 379796 54868 379848 54874
rect 379796 54810 379848 54816
rect 379520 54800 379572 54806
rect 379520 54742 379572 54748
rect 378048 54664 378100 54670
rect 378048 54606 378100 54612
rect 376024 54596 376076 54602
rect 376024 54538 376076 54544
rect 374828 54528 374880 54534
rect 374828 54470 374880 54476
rect 397472 54398 397500 57831
rect 399496 56030 399524 57831
rect 399484 56024 399536 56030
rect 399484 55966 399536 55972
rect 374644 54392 374696 54398
rect 374644 54334 374696 54340
rect 397460 54392 397512 54398
rect 397460 54334 397512 54340
rect 400232 54330 400260 57831
rect 401704 56098 401732 57831
rect 401692 56092 401744 56098
rect 401692 56034 401744 56040
rect 404372 54534 404400 57831
rect 405844 54602 405872 57831
rect 407224 55214 407252 57831
rect 408328 56574 408356 57831
rect 408316 56568 408368 56574
rect 408316 56510 408368 56516
rect 408696 56234 408724 57831
rect 408684 56228 408736 56234
rect 408684 56170 408736 56176
rect 407212 55208 407264 55214
rect 407212 55150 407264 55156
rect 409892 54670 409920 57831
rect 411258 56944 411314 56953
rect 411258 56879 411314 56888
rect 411272 56166 411300 56879
rect 411260 56160 411312 56166
rect 411260 56102 411312 56108
rect 411364 54738 411392 57831
rect 412560 56953 412588 59599
rect 416976 59566 417004 59735
rect 416964 59560 417016 59566
rect 416964 59502 417016 59508
rect 422864 59430 422892 59735
rect 423494 59664 423550 59673
rect 423494 59599 423550 59608
rect 422852 59424 422904 59430
rect 414570 59392 414626 59401
rect 414570 59327 414572 59336
rect 414624 59327 414626 59336
rect 416042 59392 416098 59401
rect 416042 59327 416098 59336
rect 418158 59392 418214 59401
rect 418158 59327 418214 59336
rect 419354 59392 419410 59401
rect 419354 59327 419410 59336
rect 420642 59392 420698 59401
rect 420642 59327 420698 59336
rect 421746 59392 421802 59401
rect 422852 59366 422904 59372
rect 421746 59327 421802 59336
rect 414572 59298 414624 59304
rect 416056 58954 416084 59327
rect 418172 59294 418200 59327
rect 418160 59288 418212 59294
rect 418160 59230 418212 59236
rect 419368 59158 419396 59327
rect 419356 59152 419408 59158
rect 419356 59094 419408 59100
rect 420656 59090 420684 59327
rect 420644 59084 420696 59090
rect 420644 59026 420696 59032
rect 421760 59022 421788 59327
rect 421748 59016 421800 59022
rect 421748 58958 421800 58964
rect 416044 58948 416096 58954
rect 416044 58890 416096 58896
rect 423508 58886 423536 59599
rect 423968 59498 423996 59735
rect 423956 59492 424008 59498
rect 423956 59434 424008 59440
rect 428186 59392 428242 59401
rect 428186 59327 428242 59336
rect 423496 58880 423548 58886
rect 423496 58822 423548 58828
rect 428200 58682 428228 59327
rect 475842 58984 475898 58993
rect 475842 58919 475898 58928
rect 468482 58848 468538 58857
rect 468482 58783 468484 58792
rect 468536 58783 468538 58792
rect 468484 58754 468536 58760
rect 475856 58750 475884 58919
rect 475844 58744 475896 58750
rect 475844 58686 475896 58692
rect 428188 58676 428240 58682
rect 428188 58618 428240 58624
rect 517624 57934 517652 165106
rect 517716 146198 517744 253166
rect 517704 146192 517756 146198
rect 517704 146134 517756 146140
rect 517808 146130 517836 253234
rect 517900 165034 517928 271186
rect 517992 253230 518020 359586
rect 519004 354674 519032 369174
rect 519096 366382 519124 400279
rect 519174 396808 519230 396817
rect 519174 396743 519230 396752
rect 519188 371958 519216 396743
rect 519358 395312 519414 395321
rect 519358 395247 519414 395256
rect 519266 394088 519322 394097
rect 519266 394023 519322 394032
rect 519176 371952 519228 371958
rect 519176 371894 519228 371900
rect 519084 366376 519136 366382
rect 519084 366318 519136 366324
rect 519280 363662 519308 394023
rect 519372 373318 519400 395247
rect 519360 373312 519412 373318
rect 519360 373254 519412 373260
rect 519372 372638 519400 373254
rect 519360 372632 519412 372638
rect 519360 372574 519412 372580
rect 519360 366376 519412 366382
rect 519360 366318 519412 366324
rect 519268 363656 519320 363662
rect 519268 363598 519320 363604
rect 518912 354646 519032 354674
rect 518912 292505 518940 354646
rect 519082 353016 519138 353025
rect 519082 352951 519138 352960
rect 518898 292496 518954 292505
rect 518898 292431 518954 292440
rect 518990 290320 519046 290329
rect 518990 290255 519046 290264
rect 517980 253224 518032 253230
rect 517980 253166 518032 253172
rect 518898 186416 518954 186425
rect 518898 186351 518954 186360
rect 517888 165028 517940 165034
rect 517888 164970 517940 164976
rect 517796 146124 517848 146130
rect 517796 146066 517848 146072
rect 517808 145586 517836 146066
rect 517796 145580 517848 145586
rect 517796 145522 517848 145528
rect 485964 57928 486016 57934
rect 415490 57896 415546 57905
rect 415490 57831 415546 57840
rect 425242 57896 425298 57905
rect 425242 57831 425298 57840
rect 426438 57896 426494 57905
rect 426438 57831 426494 57840
rect 428554 57896 428610 57905
rect 428554 57831 428610 57840
rect 429198 57896 429254 57905
rect 429198 57831 429254 57840
rect 430578 57896 430634 57905
rect 430578 57831 430634 57840
rect 432234 57896 432290 57905
rect 432234 57831 432290 57840
rect 433522 57896 433578 57905
rect 433522 57831 433578 57840
rect 434626 57896 434682 57905
rect 434626 57831 434682 57840
rect 435914 57896 435970 57905
rect 435914 57831 435970 57840
rect 436374 57896 436430 57905
rect 436374 57831 436430 57840
rect 438490 57896 438546 57905
rect 438490 57831 438546 57840
rect 445850 57896 445906 57905
rect 445850 57831 445906 57840
rect 460938 57896 460994 57905
rect 460938 57831 460994 57840
rect 465906 57896 465962 57905
rect 465906 57831 465962 57840
rect 470874 57896 470930 57905
rect 470874 57831 470876 57840
rect 415504 57254 415532 57831
rect 415492 57248 415544 57254
rect 415492 57190 415544 57196
rect 412546 56944 412602 56953
rect 412546 56879 412602 56888
rect 412638 56808 412694 56817
rect 412638 56743 412694 56752
rect 412652 56302 412680 56743
rect 412640 56296 412692 56302
rect 412640 56238 412692 56244
rect 425256 56001 425284 57831
rect 425242 55992 425298 56001
rect 425242 55927 425298 55936
rect 426452 54874 426480 57831
rect 426530 57216 426586 57225
rect 426530 57151 426586 57160
rect 426440 54868 426492 54874
rect 426440 54810 426492 54816
rect 426544 54806 426572 57151
rect 428568 56137 428596 57831
rect 428554 56128 428610 56137
rect 428554 56063 428610 56072
rect 429212 54942 429240 57831
rect 430592 55010 430620 57831
rect 430948 57316 431000 57322
rect 430948 57258 431000 57264
rect 430960 57225 430988 57258
rect 430946 57216 431002 57225
rect 430946 57151 431002 57160
rect 432248 56370 432276 57831
rect 433154 57488 433210 57497
rect 433154 57423 433210 57432
rect 433430 57488 433486 57497
rect 433536 57458 433564 57831
rect 433430 57423 433486 57432
rect 433524 57452 433576 57458
rect 433168 57225 433196 57423
rect 433154 57216 433210 57225
rect 433154 57151 433210 57160
rect 432236 56364 432288 56370
rect 432236 56306 432288 56312
rect 433444 55078 433472 57423
rect 433524 57394 433576 57400
rect 434640 56438 434668 57831
rect 434718 57488 434774 57497
rect 434718 57423 434774 57432
rect 434628 56432 434680 56438
rect 434628 56374 434680 56380
rect 433432 55072 433484 55078
rect 433432 55014 433484 55020
rect 430580 55004 430632 55010
rect 430580 54946 430632 54952
rect 429200 54936 429252 54942
rect 429200 54878 429252 54884
rect 426532 54800 426584 54806
rect 426532 54742 426584 54748
rect 411352 54732 411404 54738
rect 411352 54674 411404 54680
rect 409880 54664 409932 54670
rect 409880 54606 409932 54612
rect 405832 54596 405884 54602
rect 405832 54538 405884 54544
rect 404360 54528 404412 54534
rect 404360 54470 404412 54476
rect 434732 54466 434760 57423
rect 435928 57390 435956 57831
rect 435916 57384 435968 57390
rect 435916 57326 435968 57332
rect 436388 56506 436416 57831
rect 438504 57526 438532 57831
rect 445864 57594 445892 57831
rect 460952 57662 460980 57831
rect 465920 57730 465948 57831
rect 470928 57831 470930 57840
rect 478418 57896 478474 57905
rect 478418 57831 478474 57840
rect 485962 57896 485964 57905
rect 503260 57928 503312 57934
rect 486016 57896 486018 57905
rect 485962 57831 486018 57840
rect 503258 57896 503260 57905
rect 517612 57928 517664 57934
rect 503312 57896 503314 57905
rect 503258 57831 503314 57840
rect 503534 57896 503590 57905
rect 517612 57870 517664 57876
rect 517900 57866 517928 164970
rect 518912 79937 518940 186351
rect 519004 183433 519032 290255
rect 519096 246265 519124 352951
rect 519174 288552 519230 288561
rect 519174 288487 519230 288496
rect 519082 246256 519138 246265
rect 519082 246191 519138 246200
rect 518990 183424 519046 183433
rect 518990 183359 519046 183368
rect 518990 181928 519046 181937
rect 518990 181863 519046 181872
rect 518898 79928 518954 79937
rect 518898 79863 518954 79872
rect 519004 75449 519032 181863
rect 519096 139369 519124 246191
rect 519188 181937 519216 288487
rect 519280 287609 519308 363598
rect 519372 293865 519400 366318
rect 519464 353025 519492 459575
rect 520936 396778 520964 495450
rect 576136 405686 576164 518162
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580264 489184 580316 489190
rect 580264 489126 580316 489132
rect 580276 458153 580304 489126
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 576124 405680 576176 405686
rect 576124 405622 576176 405628
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 520924 396772 520976 396778
rect 520924 396714 520976 396720
rect 580356 396772 580408 396778
rect 580356 396714 580408 396720
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580264 378276 580316 378282
rect 580264 378218 580316 378224
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 519636 372632 519688 372638
rect 519636 372574 519688 372580
rect 519544 371952 519596 371958
rect 519544 371894 519596 371900
rect 519450 353016 519506 353025
rect 519450 352951 519506 352960
rect 519358 293856 519414 293865
rect 519358 293791 519414 293800
rect 519266 287600 519322 287609
rect 519266 287535 519322 287544
rect 519280 287094 519308 287535
rect 519268 287088 519320 287094
rect 519268 287030 519320 287036
rect 519174 181928 519230 181937
rect 519174 181863 519230 181872
rect 519280 180713 519308 287030
rect 519372 186425 519400 293791
rect 519450 292496 519506 292505
rect 519450 292431 519506 292440
rect 519358 186416 519414 186425
rect 519358 186351 519414 186360
rect 519464 184793 519492 292431
rect 519556 290329 519584 371894
rect 519542 290320 519598 290329
rect 519542 290255 519598 290264
rect 519648 288561 519676 372574
rect 580276 325281 580304 378218
rect 580368 351937 580396 396714
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 519634 288552 519690 288561
rect 519634 288487 519690 288496
rect 520186 288552 520242 288561
rect 520186 288487 520242 288496
rect 520200 288454 520228 288487
rect 520188 288448 520240 288454
rect 520188 288390 520240 288396
rect 580264 288448 580316 288454
rect 580264 288390 580316 288396
rect 580276 232393 580304 288390
rect 580356 287088 580408 287094
rect 580356 287030 580408 287036
rect 580368 272241 580396 287030
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 519450 184784 519506 184793
rect 519450 184719 519506 184728
rect 520186 184784 520242 184793
rect 520186 184719 520242 184728
rect 520200 183598 520228 184719
rect 519452 183592 519504 183598
rect 519452 183534 519504 183540
rect 520188 183592 520240 183598
rect 520188 183534 520240 183540
rect 580264 183592 580316 183598
rect 580264 183534 580316 183540
rect 519358 183424 519414 183433
rect 519358 183359 519414 183368
rect 519266 180704 519322 180713
rect 519266 180639 519322 180648
rect 519280 161474 519308 180639
rect 519188 161446 519308 161474
rect 519082 139360 519138 139369
rect 519082 139295 519138 139304
rect 518990 75440 519046 75449
rect 518990 75375 519046 75384
rect 519188 74225 519216 161446
rect 519372 76809 519400 183359
rect 519464 78305 519492 183534
rect 520096 183524 520148 183530
rect 520096 183466 520148 183472
rect 520108 183433 520136 183466
rect 520094 183424 520150 183433
rect 520094 183359 520150 183368
rect 580276 152697 580304 183534
rect 580368 183530 580396 192471
rect 580356 183524 580408 183530
rect 580356 183466 580408 183472
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580264 145648 580316 145654
rect 580264 145590 580316 145596
rect 520188 80028 520240 80034
rect 520188 79970 520240 79976
rect 520200 79937 520228 79970
rect 520186 79928 520242 79937
rect 520186 79863 520242 79872
rect 519450 78296 519506 78305
rect 519450 78231 519506 78240
rect 519358 76800 519414 76809
rect 519358 76735 519414 76744
rect 519174 74216 519230 74225
rect 519174 74151 519230 74160
rect 503534 57831 503536 57840
rect 470876 57802 470928 57808
rect 478432 57798 478460 57831
rect 503588 57831 503590 57840
rect 517888 57860 517940 57866
rect 503536 57802 503588 57808
rect 517888 57802 517940 57808
rect 478420 57792 478472 57798
rect 478420 57734 478472 57740
rect 465908 57724 465960 57730
rect 465908 57666 465960 57672
rect 460940 57656 460992 57662
rect 460940 57598 460992 57604
rect 445852 57588 445904 57594
rect 445852 57530 445904 57536
rect 438492 57520 438544 57526
rect 437478 57488 437534 57497
rect 438492 57462 438544 57468
rect 437478 57423 437534 57432
rect 436376 56500 436428 56506
rect 436376 56442 436428 56448
rect 437492 55146 437520 57423
rect 437480 55140 437532 55146
rect 437480 55082 437532 55088
rect 434720 54460 434772 54466
rect 434720 54402 434772 54408
rect 372436 54324 372488 54330
rect 372436 54266 372488 54272
rect 400220 54324 400272 54330
rect 400220 54266 400272 54272
rect 580276 33153 580304 145590
rect 580356 145580 580408 145586
rect 580356 145522 580408 145528
rect 580368 73001 580396 145522
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580460 80034 580488 112775
rect 580448 80028 580500 80034
rect 580448 79970 580500 79976
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 366364 3460 366416 3466
rect 366364 3402 366416 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 632032 3478 632088
rect 3422 579944 3478 580000
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3422 482160 3478 482216
rect 3330 410488 3386 410544
rect 3698 462576 3754 462632
rect 3606 358400 3662 358456
rect 3514 306176 3570 306232
rect 3514 97552 3570 97608
rect 3422 58520 3478 58576
rect 57610 628632 57666 628688
rect 57426 622376 57482 622432
rect 57334 597896 57390 597952
rect 57242 591776 57298 591832
rect 57150 589056 57206 589112
rect 57058 582936 57114 582992
rect 57518 619656 57574 619712
rect 57426 579672 57482 579728
rect 57794 607552 57850 607608
rect 59266 625776 59322 625832
rect 58990 616256 59046 616312
rect 57886 604016 57942 604072
rect 57794 595176 57850 595232
rect 57794 573416 57850 573472
rect 58898 601296 58954 601352
rect 58530 576816 58586 576872
rect 58806 585656 58862 585712
rect 59174 613536 59230 613592
rect 59082 610136 59138 610192
rect 59542 570732 59598 570788
rect 68098 552608 68154 552664
rect 120814 606328 120870 606384
rect 121090 591164 121146 591220
rect 121182 578924 121238 578980
rect 121550 570016 121606 570072
rect 121826 621152 121882 621208
rect 121734 615576 121790 615632
rect 121918 608912 121974 608968
rect 122010 593952 122066 594008
rect 122102 587968 122158 588024
rect 122838 627952 122894 628008
rect 122286 572736 122342 572792
rect 123022 625232 123078 625288
rect 123114 612720 123170 612776
rect 123298 603064 123354 603120
rect 123206 600344 123262 600400
rect 124126 596672 124182 596728
rect 123390 584432 123446 584488
rect 123482 581712 123538 581768
rect 123482 575592 123538 575648
rect 146298 628632 146354 628688
rect 147310 622376 147366 622432
rect 146298 619676 146354 619712
rect 146298 619656 146300 619676
rect 146300 619656 146352 619676
rect 146352 619656 146354 619676
rect 146298 616256 146354 616312
rect 146850 613536 146906 613592
rect 146206 604152 146262 604208
rect 146298 597896 146354 597952
rect 146298 585656 146354 585712
rect 146298 582936 146354 582992
rect 146298 579692 146354 579728
rect 146298 579672 146300 579692
rect 146300 579672 146352 579692
rect 146352 579672 146354 579692
rect 147126 595176 147182 595232
rect 147034 576816 147090 576872
rect 147218 589056 147274 589112
rect 147586 607552 147642 607608
rect 148230 570696 148286 570752
rect 148690 625776 148746 625832
rect 148506 610136 148562 610192
rect 148414 591776 148470 591832
rect 148598 601296 148654 601352
rect 149058 573416 149114 573472
rect 211250 627952 211306 628008
rect 211158 615576 211214 615632
rect 210790 575592 210846 575648
rect 210882 570288 210938 570344
rect 211434 618432 211490 618488
rect 211342 612720 211398 612776
rect 211618 606328 211674 606384
rect 211526 600344 211582 600400
rect 211710 593952 211766 594008
rect 211802 584432 211858 584488
rect 212538 581712 212594 581768
rect 212722 625232 212778 625288
rect 213274 621152 213330 621208
rect 212814 608912 212870 608968
rect 212906 603064 212962 603120
rect 213090 590688 213146 590744
rect 212998 587968 213054 588024
rect 213182 578312 213238 578368
rect 213366 572736 213422 572792
rect 214102 596672 214158 596728
rect 237378 628632 237434 628688
rect 237378 622412 237380 622432
rect 237380 622412 237432 622432
rect 237432 622412 237434 622432
rect 237378 622376 237434 622412
rect 237378 619676 237434 619712
rect 237378 619656 237380 619676
rect 237380 619656 237432 619676
rect 237432 619656 237434 619676
rect 237378 616256 237434 616312
rect 237378 613536 237434 613592
rect 237378 610136 237434 610192
rect 238022 604152 238078 604208
rect 237378 601296 237434 601352
rect 237378 597896 237434 597952
rect 237378 595176 237434 595232
rect 237378 591776 237434 591832
rect 237378 589056 237434 589112
rect 237378 585656 237434 585712
rect 236734 582936 236790 582992
rect 237378 579692 237434 579728
rect 237378 579672 237380 579692
rect 237380 579672 237432 579692
rect 237432 579672 237434 579692
rect 237378 576852 237380 576872
rect 237380 576852 237432 576872
rect 237432 576852 237434 576872
rect 237378 576816 237434 576852
rect 237378 573416 237434 573472
rect 237378 570696 237434 570752
rect 237194 548120 237250 548176
rect 238298 625776 238354 625832
rect 238942 607552 238998 607608
rect 300858 628088 300914 628144
rect 238666 549480 238722 549536
rect 241518 549616 241574 549672
rect 245842 549888 245898 549944
rect 248694 549752 248750 549808
rect 255134 549344 255190 549400
rect 300950 625368 301006 625424
rect 302882 621152 302938 621208
rect 301134 618432 301190 618488
rect 301042 615576 301098 615632
rect 301226 612720 301282 612776
rect 302422 608912 302478 608968
rect 301318 600344 301374 600400
rect 301410 593952 301466 594008
rect 302238 587968 302294 588024
rect 301502 581712 301558 581768
rect 301594 575592 301650 575648
rect 301686 570016 301742 570072
rect 302330 578312 302386 578368
rect 302514 603064 302570 603120
rect 302698 596672 302754 596728
rect 302606 590688 302662 590744
rect 302790 584432 302846 584488
rect 293774 548120 293830 548176
rect 298098 550160 298154 550216
rect 297362 550024 297418 550080
rect 301502 520104 301558 520160
rect 301778 549752 301834 549808
rect 301962 549616 302018 549672
rect 301870 547848 301926 547904
rect 302606 540368 302662 540424
rect 301962 522416 302018 522472
rect 57886 517928 57942 517984
rect 43902 482296 43958 482352
rect 42614 479984 42670 480040
rect 43718 477128 43774 477184
rect 43534 476856 43590 476912
rect 43626 476720 43682 476776
rect 43810 476992 43866 477048
rect 43994 378800 44050 378856
rect 46570 482568 46626 482624
rect 46478 482432 46534 482488
rect 46018 272448 46074 272504
rect 46570 270952 46626 271008
rect 47582 380024 47638 380080
rect 47766 379344 47822 379400
rect 47674 379208 47730 379264
rect 47582 378936 47638 378992
rect 47766 378936 47822 378992
rect 47674 271496 47730 271552
rect 47858 271360 47914 271416
rect 49054 271632 49110 271688
rect 49238 165416 49294 165472
rect 49514 471144 49570 471200
rect 49330 165280 49386 165336
rect 49514 165144 49570 165200
rect 50158 272992 50214 273048
rect 50250 272856 50306 272912
rect 50986 380704 51042 380760
rect 50986 379480 51042 379536
rect 50250 145560 50306 145616
rect 51630 271768 51686 271824
rect 51998 465160 52054 465216
rect 302974 606328 303030 606384
rect 303066 572736 303122 572792
rect 302974 525408 303030 525464
rect 302698 510448 302754 510504
rect 302238 495508 302294 495544
rect 302238 495488 302240 495508
rect 302240 495488 302292 495508
rect 302292 495488 302294 495508
rect 53286 484472 53342 484528
rect 53654 484472 53710 484528
rect 52366 388456 52422 388512
rect 52458 272720 52514 272776
rect 53010 271768 53066 271824
rect 53286 270408 53342 270464
rect 54390 375400 54446 375456
rect 54206 282240 54262 282296
rect 53838 271088 53894 271144
rect 54390 271088 54446 271144
rect 55126 471552 55182 471608
rect 54482 145832 54538 145888
rect 54574 145560 54630 145616
rect 55678 465160 55734 465216
rect 56138 471280 56194 471336
rect 56966 417152 57022 417208
rect 57058 391448 57114 391504
rect 57058 389036 57060 389056
rect 57060 389036 57112 389056
rect 57112 389036 57114 389056
rect 57058 389000 57114 389036
rect 56874 309032 56930 309088
rect 56874 307808 56930 307864
rect 56782 307672 56838 307728
rect 56782 203496 56838 203552
rect 56230 146240 56286 146296
rect 56322 145696 56378 145752
rect 56874 201320 56930 201376
rect 57518 389272 57574 389328
rect 57518 311072 57574 311128
rect 57334 310392 57390 310448
rect 57242 282512 57298 282568
rect 57242 268912 57298 268968
rect 57150 204176 57206 204232
rect 57058 195200 57114 195256
rect 56782 96464 56838 96520
rect 57426 301552 57482 301608
rect 57334 203496 57390 203552
rect 57334 198736 57390 198792
rect 57150 97416 57206 97472
rect 57886 417288 57942 417344
rect 57886 414160 57942 414216
rect 57886 413208 57942 413264
rect 57886 411440 57942 411496
rect 57886 410352 57942 410408
rect 57886 408584 57942 408640
rect 58622 388456 58678 388512
rect 57794 310392 57850 310448
rect 57702 309032 57758 309088
rect 57794 307672 57850 307728
rect 57794 306720 57850 306776
rect 57702 304952 57758 305008
rect 57610 303612 57666 303648
rect 57610 303592 57612 303612
rect 57612 303592 57664 303612
rect 57664 303592 57666 303612
rect 57518 204176 57574 204232
rect 57610 201320 57666 201376
rect 57426 196288 57482 196344
rect 57334 93336 57390 93392
rect 57518 164092 57520 164112
rect 57520 164092 57572 164112
rect 57572 164092 57574 164112
rect 57518 164056 57574 164092
rect 57886 282512 57942 282568
rect 57794 199824 57850 199880
rect 57794 198736 57850 198792
rect 57794 198056 57850 198112
rect 57702 195200 57758 195256
rect 57610 93744 57666 93800
rect 57426 90480 57482 90536
rect 58714 284144 58770 284200
rect 58806 281968 58862 282024
rect 57886 175752 57942 175808
rect 57794 91024 57850 91080
rect 57702 88168 57758 88224
rect 57610 70080 57666 70136
rect 58714 147736 58770 147792
rect 58898 177520 58954 177576
rect 58806 146240 58862 146296
rect 57886 68856 57942 68912
rect 3422 19352 3478 19408
rect 58990 145832 59046 145888
rect 59818 471688 59874 471744
rect 59450 272584 59506 272640
rect 59358 269048 59414 269104
rect 59450 175888 59506 175944
rect 62210 478080 62266 478136
rect 66350 482840 66406 482896
rect 66258 466384 66314 466440
rect 68926 484880 68982 484936
rect 67822 469784 67878 469840
rect 67730 469104 67786 469160
rect 69018 465840 69074 465896
rect 69202 468968 69258 469024
rect 72514 485696 72570 485752
rect 71870 467064 71926 467120
rect 71778 466248 71834 466304
rect 73802 485560 73858 485616
rect 74262 485424 74318 485480
rect 74446 485424 74502 485480
rect 73158 467200 73214 467256
rect 74538 466112 74594 466168
rect 76010 485288 76066 485344
rect 77298 485152 77354 485208
rect 78678 468832 78734 468888
rect 78770 468696 78826 468752
rect 79966 485424 80022 485480
rect 80518 479984 80574 480040
rect 78862 468560 78918 468616
rect 80242 468424 80298 468480
rect 81530 471416 81586 471472
rect 88430 471552 88486 471608
rect 89810 471280 89866 471336
rect 91374 485016 91430 485072
rect 76010 465976 76066 466032
rect 74630 465704 74686 465760
rect 69110 465568 69166 465624
rect 92662 471688 92718 471744
rect 94226 471144 94282 471200
rect 118790 479848 118846 479904
rect 117962 479576 118018 479632
rect 120446 482704 120502 482760
rect 120906 482568 120962 482624
rect 120078 482432 120134 482488
rect 121366 482296 121422 482352
rect 118882 479440 118938 479496
rect 122378 479712 122434 479768
rect 124310 477128 124366 477184
rect 125690 476992 125746 477048
rect 125782 476856 125838 476912
rect 127070 476720 127126 476776
rect 125598 464344 125654 464400
rect 145654 485288 145710 485344
rect 145470 485016 145526 485072
rect 147586 485152 147642 485208
rect 147218 480800 147274 480856
rect 145746 476856 145802 476912
rect 143630 474000 143686 474056
rect 143538 472504 143594 472560
rect 150254 483656 150310 483712
rect 147770 479576 147826 479632
rect 151358 476720 151414 476776
rect 150438 475360 150494 475416
rect 147678 469784 147734 469840
rect 152738 478216 152794 478272
rect 156510 483792 156566 483848
rect 155866 482296 155922 482352
rect 155222 480936 155278 480992
rect 154026 479440 154082 479496
rect 158626 485696 158682 485752
rect 157522 475496 157578 475552
rect 161570 471280 161626 471336
rect 161478 468424 161534 468480
rect 155958 467064 156014 467120
rect 163686 485424 163742 485480
rect 162858 465840 162914 465896
rect 165802 466112 165858 466168
rect 167090 468832 167146 468888
rect 169850 472640 169906 472696
rect 171138 485560 171194 485616
rect 169942 471688 169998 471744
rect 169758 471552 169814 471608
rect 171230 472776 171286 472832
rect 171138 471144 171194 471200
rect 172518 468968 172574 469024
rect 168562 468696 168618 468752
rect 168378 468560 168434 468616
rect 166998 465976 167054 466032
rect 174818 471416 174874 471472
rect 178682 479712 178738 479768
rect 180154 467236 180156 467256
rect 180156 467236 180208 467256
rect 180208 467236 180210 467256
rect 180154 467200 180210 467236
rect 178038 466540 178094 466576
rect 178038 466520 178040 466540
rect 178040 466520 178092 466540
rect 178092 466520 178094 466540
rect 182270 485696 182326 485752
rect 182822 466248 182878 466304
rect 165618 465704 165674 465760
rect 184846 485696 184902 485752
rect 187054 484880 187110 484936
rect 191102 485152 191158 485208
rect 191102 484608 191158 484664
rect 190918 466520 190974 466576
rect 60002 380976 60058 381032
rect 59450 140800 59506 140856
rect 93398 380840 93454 380896
rect 110970 380840 111026 380896
rect 113546 380840 113602 380896
rect 116030 380840 116086 380896
rect 118422 380840 118478 380896
rect 120998 380840 121054 380896
rect 123482 380840 123538 380896
rect 125966 380840 126022 380896
rect 131026 380840 131082 380896
rect 133510 380840 133566 380896
rect 135902 380840 135958 380896
rect 143538 380876 143540 380896
rect 143540 380876 143592 380896
rect 143592 380876 143594 380896
rect 143538 380840 143594 380876
rect 146022 380840 146078 380896
rect 158534 380840 158590 380896
rect 160926 380840 160982 380896
rect 163410 380840 163466 380896
rect 165986 380840 166042 380896
rect 85486 379344 85542 379400
rect 86590 379344 86646 379400
rect 87694 379344 87750 379400
rect 88338 379364 88394 379400
rect 88338 379344 88340 379364
rect 88340 379344 88392 379364
rect 88392 379344 88394 379364
rect 80426 379208 80482 379264
rect 81438 379208 81494 379264
rect 80426 378392 80482 378448
rect 83462 378800 83518 378856
rect 88798 379364 88854 379400
rect 88798 379344 88800 379364
rect 88800 379344 88852 379364
rect 88852 379344 88854 379364
rect 90086 379344 90142 379400
rect 90638 379344 90694 379400
rect 91374 379344 91430 379400
rect 92386 379344 92442 379400
rect 128358 380296 128414 380352
rect 155958 380296 156014 380352
rect 93490 379380 93492 379400
rect 93492 379380 93544 379400
rect 93544 379380 93546 379400
rect 93490 379344 93546 379380
rect 96066 379344 96122 379400
rect 98274 379344 98330 379400
rect 98458 379344 98514 379400
rect 101034 379344 101090 379400
rect 103518 379344 103574 379400
rect 105266 379344 105322 379400
rect 108210 379344 108266 379400
rect 108854 379344 108910 379400
rect 111246 379344 111302 379400
rect 112626 379344 112682 379400
rect 113454 379344 113510 379400
rect 114466 379344 114522 379400
rect 117134 379344 117190 379400
rect 141054 379344 141110 379400
rect 148598 379344 148654 379400
rect 150990 379344 151046 379400
rect 153566 379344 153622 379400
rect 183190 379344 183246 379400
rect 95974 379208 96030 379264
rect 94686 378664 94742 378720
rect 85026 378120 85082 378176
rect 97170 378664 97226 378720
rect 99470 379208 99526 379264
rect 102966 379208 103022 379264
rect 101862 378120 101918 378176
rect 105542 379208 105598 379264
rect 104438 378256 104494 378312
rect 138478 378664 138534 378720
rect 107566 378256 107622 378312
rect 106462 378120 106518 378176
rect 182270 378120 182326 378176
rect 182822 378120 182878 378176
rect 178682 358808 178738 358864
rect 179878 358808 179934 358864
rect 197358 485188 197360 485208
rect 197360 485188 197412 485208
rect 197412 485188 197414 485208
rect 197358 485152 197414 485188
rect 197358 484744 197414 484800
rect 190918 358808 190974 358864
rect 95974 273808 96030 273864
rect 113362 273808 113418 273864
rect 76010 273128 76066 273184
rect 77114 273128 77170 273184
rect 90730 273128 90786 273184
rect 93674 273128 93730 273184
rect 94226 273128 94282 273184
rect 94226 272856 94282 272912
rect 94410 272856 94466 272912
rect 95882 272856 95938 272912
rect 83002 272332 83058 272368
rect 83002 272312 83004 272332
rect 83004 272312 83056 272332
rect 83056 272312 83058 272332
rect 98458 272856 98514 272912
rect 100758 272312 100814 272368
rect 99378 272176 99434 272232
rect 84198 271768 84254 271824
rect 97998 271768 98054 271824
rect 62118 271088 62174 271144
rect 88338 270972 88394 271008
rect 88338 270952 88340 270972
rect 88340 270952 88392 270972
rect 88392 270952 88394 270972
rect 89718 270952 89774 271008
rect 85578 270816 85634 270872
rect 88338 270816 88394 270872
rect 84658 270544 84714 270600
rect 86958 270544 87014 270600
rect 92478 270816 92534 270872
rect 91098 270544 91154 270600
rect 102138 271768 102194 271824
rect 104898 271768 104954 271824
rect 107474 271768 107530 271824
rect 100758 271632 100814 271688
rect 110418 271632 110474 271688
rect 103518 271360 103574 271416
rect 113178 271380 113234 271416
rect 113178 271360 113180 271380
rect 113180 271360 113232 271380
rect 113232 271360 113234 271380
rect 104898 271224 104954 271280
rect 107658 271244 107714 271280
rect 107658 271224 107660 271244
rect 107660 271224 107712 271244
rect 107712 271224 107714 271244
rect 111798 271088 111854 271144
rect 106278 270816 106334 270872
rect 109038 270544 109094 270600
rect 110418 270544 110474 270600
rect 133418 273672 133474 273728
rect 135902 273556 135958 273592
rect 135902 273536 135904 273556
rect 135904 273536 135956 273556
rect 135956 273536 135958 273556
rect 138478 273536 138534 273592
rect 140870 273536 140926 273592
rect 143538 273536 143594 273592
rect 145930 273536 145986 273592
rect 114466 271768 114522 271824
rect 123206 271788 123262 271824
rect 123206 271768 123208 271788
rect 123208 271768 123260 271788
rect 123260 271768 123262 271788
rect 125598 271768 125654 271824
rect 120078 271632 120134 271688
rect 115938 271516 115994 271552
rect 115938 271496 115940 271516
rect 115940 271496 115992 271516
rect 115992 271496 115994 271516
rect 117318 271496 117374 271552
rect 118698 271224 118754 271280
rect 114558 270952 114614 271008
rect 115938 270816 115994 270872
rect 129738 271804 129740 271824
rect 129740 271804 129792 271824
rect 129792 271804 129794 271824
rect 129738 271768 129794 271804
rect 151358 271768 151414 271824
rect 154486 271804 154488 271824
rect 154488 271804 154540 271824
rect 154540 271804 154542 271824
rect 154486 271768 154542 271804
rect 158626 271788 158682 271824
rect 158626 271768 158628 271788
rect 158628 271768 158680 271788
rect 158680 271768 158682 271788
rect 128358 271652 128414 271688
rect 128358 271632 128360 271652
rect 128360 271632 128412 271652
rect 128412 271632 128414 271652
rect 157246 271652 157302 271688
rect 157246 271632 157248 271652
rect 157248 271632 157300 271652
rect 157300 271632 157302 271652
rect 161294 271632 161350 271688
rect 164146 271632 164202 271688
rect 166906 271632 166962 271688
rect 183466 271632 183522 271688
rect 147678 270816 147734 270872
rect 183466 270564 183522 270600
rect 183466 270544 183468 270564
rect 183468 270544 183520 270564
rect 183520 270544 183522 270564
rect 180154 253308 180156 253328
rect 180156 253308 180208 253328
rect 180208 253308 180210 253328
rect 180154 253272 180210 253308
rect 179326 253136 179382 253192
rect 191746 253172 191748 253192
rect 191748 253172 191800 253192
rect 191800 253172 191802 253192
rect 191746 253136 191802 253172
rect 96066 166776 96122 166832
rect 98458 166776 98514 166832
rect 101034 166812 101036 166832
rect 101036 166812 101088 166832
rect 101088 166812 101090 166832
rect 101034 166776 101090 166812
rect 105818 166796 105874 166832
rect 105818 166776 105820 166796
rect 105820 166776 105872 166796
rect 105872 166776 105874 166796
rect 108210 166776 108266 166832
rect 138478 166776 138534 166832
rect 140870 166776 140926 166832
rect 145930 166776 145986 166832
rect 111154 166504 111210 166560
rect 116950 166504 117006 166560
rect 163318 166640 163374 166696
rect 148506 166504 148562 166560
rect 153290 166388 153346 166424
rect 153290 166368 153292 166388
rect 153292 166368 153344 166388
rect 153344 166368 153346 166388
rect 81438 165552 81494 165608
rect 84198 165552 84254 165608
rect 91190 165552 91246 165608
rect 95238 165552 95294 165608
rect 99378 165552 99434 165608
rect 103518 165552 103574 165608
rect 109314 165552 109370 165608
rect 110970 165552 111026 165608
rect 113546 165552 113602 165608
rect 115938 165552 115994 165608
rect 117870 165552 117926 165608
rect 118146 165552 118202 165608
rect 120906 165552 120962 165608
rect 123482 165552 123538 165608
rect 125874 165552 125930 165608
rect 128358 165552 128414 165608
rect 129738 165552 129794 165608
rect 132498 165552 132554 165608
rect 135258 165552 135314 165608
rect 150438 165572 150494 165608
rect 150438 165552 150440 165572
rect 150440 165552 150492 165572
rect 150492 165552 150494 165572
rect 75918 164328 75974 164384
rect 76010 164192 76066 164248
rect 77298 164192 77354 164248
rect 78678 164192 78734 164248
rect 80058 164192 80114 164248
rect 82818 164192 82874 164248
rect 88338 164736 88394 164792
rect 89994 164756 90050 164792
rect 89994 164736 89996 164756
rect 89996 164736 90048 164756
rect 90048 164736 90050 164756
rect 84290 164192 84346 164248
rect 85578 164192 85634 164248
rect 86958 164192 87014 164248
rect 88430 164192 88486 164248
rect 89810 164192 89866 164248
rect 91098 164192 91154 164248
rect 92478 164192 92534 164248
rect 93858 164192 93914 164248
rect 96618 164464 96674 164520
rect 97998 164192 98054 164248
rect 100758 164348 100814 164384
rect 100758 164328 100760 164348
rect 100760 164328 100812 164348
rect 100812 164328 100814 164348
rect 103518 164328 103574 164384
rect 100758 164192 100814 164248
rect 102138 164192 102194 164248
rect 106186 164192 106242 164248
rect 106370 164192 106426 164248
rect 107566 164192 107622 164248
rect 107658 164056 107714 164112
rect 114466 164892 114522 164928
rect 114466 164872 114468 164892
rect 114468 164872 114520 164892
rect 114520 164872 114522 164892
rect 112074 164600 112130 164656
rect 114650 164464 114706 164520
rect 115754 164600 115810 164656
rect 183190 165552 183246 165608
rect 183466 165552 183522 165608
rect 118882 165008 118938 165064
rect 102138 146240 102194 146296
rect 100758 145832 100814 145888
rect 99378 145696 99434 145752
rect 98642 145560 98698 145616
rect 179050 144880 179106 144936
rect 179694 144880 179750 144936
rect 191286 144880 191342 144936
rect 77114 59764 77170 59800
rect 77114 59744 77116 59764
rect 77116 59744 77168 59764
rect 77168 59744 77170 59764
rect 83094 59744 83150 59800
rect 101770 59744 101826 59800
rect 103886 59744 103942 59800
rect 107566 59744 107622 59800
rect 113546 59744 113602 59800
rect 94502 59608 94558 59664
rect 96986 59608 97042 59664
rect 98090 59608 98146 59664
rect 100758 59628 100814 59664
rect 100758 59608 100760 59628
rect 100760 59608 100812 59628
rect 100812 59608 100814 59628
rect 95882 59472 95938 59528
rect 102782 59608 102838 59664
rect 108670 59608 108726 59664
rect 110970 59336 111026 59392
rect 148506 59200 148562 59256
rect 150898 59200 150954 59256
rect 84198 57976 84254 58032
rect 76010 57840 76066 57896
rect 78218 57840 78274 57896
rect 79506 57840 79562 57896
rect 80058 57840 80114 57896
rect 81898 57840 81954 57896
rect 85394 57840 85450 57896
rect 86498 57840 86554 57896
rect 86958 57840 87014 57896
rect 88706 57840 88762 57896
rect 89810 57840 89866 57896
rect 90730 57840 90786 57896
rect 91190 57840 91246 57896
rect 92202 57840 92258 57896
rect 92478 57840 92534 57896
rect 93582 57840 93638 57896
rect 99378 57840 99434 57896
rect 109498 57840 109554 57896
rect 112074 57840 112130 57896
rect 113822 57840 113878 57896
rect 115938 57840 115994 57896
rect 116674 57840 116730 57896
rect 123482 57840 123538 57896
rect 125874 57840 125930 57896
rect 128358 57840 128414 57896
rect 130842 57840 130898 57896
rect 133418 57840 133474 57896
rect 145562 57860 145618 57896
rect 145562 57840 145564 57860
rect 145564 57840 145616 57860
rect 145616 57840 145618 57860
rect 98550 57432 98606 57488
rect 106278 57568 106334 57624
rect 98550 57160 98606 57216
rect 110418 57568 110474 57624
rect 113270 57568 113326 57624
rect 114558 57568 114614 57624
rect 118698 57568 118754 57624
rect 153290 57840 153346 57896
rect 183282 57860 183338 57896
rect 183282 57840 183284 57860
rect 183284 57840 183336 57860
rect 183336 57840 183338 57860
rect 198186 397976 198242 398032
rect 198922 460128 198978 460184
rect 199198 398112 199254 398168
rect 199106 396752 199162 396808
rect 199014 379344 199070 379400
rect 199198 396072 199254 396128
rect 200210 485288 200266 485344
rect 200486 484744 200542 484800
rect 199566 400288 199622 400344
rect 199474 377848 199530 377904
rect 199382 371864 199438 371920
rect 198830 353096 198886 353152
rect 198738 290944 198794 291000
rect 198922 291624 198978 291680
rect 198830 246200 198886 246256
rect 198738 183504 198794 183560
rect 198738 182008 198794 182064
rect 199198 292712 199254 292768
rect 199014 288768 199070 288824
rect 198922 184864 198978 184920
rect 198922 183504 198978 183560
rect 198830 139168 198886 139224
rect 199106 288360 199162 288416
rect 199106 287544 199162 287600
rect 199014 182008 199070 182064
rect 199750 394576 199806 394632
rect 199474 291624 199530 291680
rect 199658 292712 199714 292768
rect 199750 290944 199806 291000
rect 199566 288360 199622 288416
rect 201498 484916 201500 484936
rect 201500 484916 201552 484936
rect 201552 484916 201554 484936
rect 201498 484880 201554 484916
rect 199290 186360 199346 186416
rect 199198 184864 199254 184920
rect 199106 180648 199162 180704
rect 198922 76336 198978 76392
rect 198738 74840 198794 74896
rect 202786 379480 202842 379536
rect 199290 79328 199346 79384
rect 199198 77696 199254 77752
rect 199014 73616 199070 73672
rect 203062 380296 203118 380352
rect 204442 485152 204498 485208
rect 204350 380568 204406 380624
rect 204902 471280 204958 471336
rect 204994 466112 205050 466168
rect 205546 411304 205602 411360
rect 206190 485152 206246 485208
rect 206190 380976 206246 381032
rect 206466 465976 206522 466032
rect 206834 378528 206890 378584
rect 207570 379072 207626 379128
rect 207570 270272 207626 270328
rect 207938 379072 207994 379128
rect 207938 378800 207994 378856
rect 208122 380160 208178 380216
rect 208398 485052 208400 485072
rect 208400 485052 208452 485072
rect 208452 485052 208454 485072
rect 208398 485016 208454 485052
rect 208398 484780 208400 484800
rect 208400 484780 208452 484800
rect 208452 484780 208454 484800
rect 208398 484744 208454 484780
rect 208674 390632 208730 390688
rect 208214 378664 208270 378720
rect 207754 270952 207810 271008
rect 208306 270272 208362 270328
rect 183466 57740 183468 57760
rect 183468 57740 183520 57760
rect 183520 57740 183522 57760
rect 183466 57704 183522 57740
rect 208858 378936 208914 378992
rect 208858 269728 208914 269784
rect 209594 379480 209650 379536
rect 209502 375400 209558 375456
rect 211158 485732 211160 485752
rect 211160 485732 211212 485752
rect 211212 485732 211214 485752
rect 211158 485696 211214 485732
rect 209962 469104 210018 469160
rect 211158 484608 211214 484664
rect 155958 57568 156014 57624
rect 160098 57568 160154 57624
rect 165618 57568 165674 57624
rect 153290 56208 153346 56264
rect 212538 485560 212594 485616
rect 210974 375536 211030 375592
rect 210882 270136 210938 270192
rect 211066 375400 211122 375456
rect 211710 379072 211766 379128
rect 211526 270408 211582 270464
rect 211986 468696 212042 468752
rect 212078 271632 212134 271688
rect 212814 380296 212870 380352
rect 212630 378528 212686 378584
rect 212446 378120 212502 378176
rect 212630 378120 212686 378176
rect 212354 269728 212410 269784
rect 212630 376388 212632 376408
rect 212632 376388 212684 376408
rect 212684 376388 212686 376408
rect 212630 376352 212686 376388
rect 212814 271768 212870 271824
rect 213734 380296 213790 380352
rect 213366 271768 213422 271824
rect 213366 271360 213422 271416
rect 213550 376388 213552 376408
rect 213552 376388 213604 376408
rect 213604 376388 213606 376408
rect 213550 376352 213606 376388
rect 165618 55120 165674 55176
rect 160098 54984 160154 55040
rect 155958 54848 156014 54904
rect 118698 54712 118754 54768
rect 213826 379208 213882 379264
rect 213826 378256 213882 378312
rect 214746 484472 214802 484528
rect 213826 376760 213882 376816
rect 213458 145560 213514 145616
rect 214194 146240 214250 146296
rect 215114 375536 215170 375592
rect 214930 270136 214986 270192
rect 213734 55120 213790 55176
rect 214930 146240 214986 146296
rect 215206 375400 215262 375456
rect 215482 380840 215538 380896
rect 215666 273264 215722 273320
rect 216126 465840 216182 465896
rect 216678 417832 216734 417888
rect 217138 414704 217194 414760
rect 216862 413752 216918 413808
rect 216770 410896 216826 410952
rect 216678 390904 216734 390960
rect 216678 389272 216734 389328
rect 216678 389000 216734 389056
rect 216586 380840 216642 380896
rect 216678 380704 216734 380760
rect 216678 379616 216734 379672
rect 217230 411304 217286 411360
rect 217322 409128 217378 409184
rect 217138 380024 217194 380080
rect 217138 379480 217194 379536
rect 217138 309984 217194 310040
rect 217046 307672 217102 307728
rect 216770 304952 216826 305008
rect 216678 284008 216734 284064
rect 216678 282240 216734 282296
rect 216954 302096 217010 302152
rect 216862 282104 216918 282160
rect 216770 198056 216826 198112
rect 216770 196968 216826 197024
rect 216678 176976 216734 177032
rect 216678 175344 216734 175400
rect 216586 145968 216642 146024
rect 214930 54984 214986 55040
rect 216954 195200 217010 195256
rect 216954 175072 217010 175128
rect 217414 377848 217470 377904
rect 217322 304952 217378 305008
rect 217230 268640 217286 268696
rect 217690 411984 217746 412040
rect 217690 411304 217746 411360
rect 217966 416880 218022 416936
rect 217874 409128 217930 409184
rect 217874 379616 217930 379672
rect 217690 379480 217746 379536
rect 217506 374856 217562 374912
rect 217506 310936 217562 310992
rect 217506 307672 217562 307728
rect 217506 306720 217562 306776
rect 217414 203904 217470 203960
rect 217138 202952 217194 203008
rect 217230 198736 217286 198792
rect 216770 89936 216826 89992
rect 216678 69944 216734 70000
rect 216678 68312 216734 68368
rect 217322 162596 217324 162616
rect 217324 162596 217376 162616
rect 217376 162596 217378 162616
rect 217322 162560 217378 162596
rect 217690 307808 217746 307864
rect 217598 203904 217654 203960
rect 217598 202952 217654 203008
rect 217506 199824 217562 199880
rect 217506 198736 217562 198792
rect 217506 198056 217562 198112
rect 217414 96872 217470 96928
rect 217230 92792 217286 92848
rect 217782 303864 217838 303920
rect 217690 200776 217746 200832
rect 217598 95920 217654 95976
rect 218334 379072 218390 379128
rect 218334 378528 218390 378584
rect 217966 309984 218022 310040
rect 217782 196968 217838 197024
rect 217782 195200 217838 195256
rect 217690 93744 217746 93800
rect 217506 91024 217562 91080
rect 217782 88168 217838 88224
rect 218242 165552 218298 165608
rect 217966 68312 218022 68368
rect 218610 146104 218666 146160
rect 218978 465704 219034 465760
rect 219070 269884 219126 269920
rect 219070 269864 219072 269884
rect 219072 269864 219124 269884
rect 219124 269864 219126 269884
rect 219070 60560 219126 60616
rect 219898 145832 219954 145888
rect 222566 482296 222622 482352
rect 225694 485152 225750 485208
rect 226154 485016 226210 485072
rect 224866 484472 224922 484528
rect 223670 478216 223726 478272
rect 223578 474000 223634 474056
rect 227994 476856 228050 476912
rect 227718 474408 227774 474464
rect 230662 485560 230718 485616
rect 230386 483656 230442 483712
rect 231766 485016 231822 485072
rect 232318 485152 232374 485208
rect 232134 480800 232190 480856
rect 234342 485424 234398 485480
rect 233330 479576 233386 479632
rect 235814 485696 235870 485752
rect 235906 485288 235962 485344
rect 234618 476720 234674 476776
rect 230754 474136 230810 474192
rect 229098 472504 229154 472560
rect 236366 482432 236422 482488
rect 240230 474272 240286 474328
rect 247314 480936 247370 480992
rect 248694 484880 248750 484936
rect 252926 483792 252982 483848
rect 256330 475360 256386 475416
rect 265070 468424 265126 468480
rect 276110 474544 276166 474600
rect 281078 483928 281134 483984
rect 292578 467064 292634 467120
rect 294142 475496 294198 475552
rect 297178 476992 297234 477048
rect 317234 547984 317290 548040
rect 320822 550568 320878 550624
rect 321098 632168 321154 632224
rect 321558 627408 321614 627464
rect 321558 622648 321614 622704
rect 321558 617888 321614 617944
rect 321558 613128 321614 613184
rect 321558 608368 321614 608424
rect 321558 603608 321614 603664
rect 321558 598848 321614 598904
rect 321558 589348 321614 589384
rect 321558 589328 321560 589348
rect 321560 589328 321612 589348
rect 321612 589328 321614 589348
rect 321558 584568 321614 584624
rect 321558 579808 321614 579864
rect 321558 574368 321614 574424
rect 321558 569608 321614 569664
rect 321558 564848 321614 564904
rect 321558 560088 321614 560144
rect 321558 555328 321614 555384
rect 320914 550160 320970 550216
rect 322202 550024 322258 550080
rect 321098 549344 321154 549400
rect 321834 545808 321890 545864
rect 321558 541048 321614 541104
rect 321558 536288 321614 536344
rect 322202 531528 322258 531584
rect 321558 526768 321614 526824
rect 324778 634888 324834 634944
rect 324226 594088 324282 594144
rect 423862 634888 423918 634944
rect 333058 632576 333114 632632
rect 351090 632440 351146 632496
rect 433338 619112 433394 619168
rect 433338 589464 433394 589520
rect 323674 549888 323730 549944
rect 329746 519968 329802 520024
rect 316682 482160 316738 482216
rect 338486 466520 338542 466576
rect 339774 466540 339830 466576
rect 339774 466520 339776 466540
rect 339776 466520 339828 466540
rect 339828 466520 339830 466540
rect 350998 466520 351054 466576
rect 235998 380704 236054 380760
rect 237102 380704 237158 380760
rect 243082 380704 243138 380760
rect 245382 380704 245438 380760
rect 256054 380704 256110 380760
rect 269762 380704 269818 380760
rect 221094 378392 221150 378448
rect 254490 380568 254546 380624
rect 255870 380568 255926 380624
rect 256974 380568 257030 380624
rect 259458 380568 259514 380624
rect 265254 380568 265310 380624
rect 246026 379344 246082 379400
rect 247498 379344 247554 379400
rect 248602 379344 248658 379400
rect 250074 379344 250130 379400
rect 251178 379344 251234 379400
rect 252282 379344 252338 379400
rect 253386 379344 253442 379400
rect 258078 379344 258134 379400
rect 261666 379344 261722 379400
rect 248234 378800 248290 378856
rect 244278 378256 244334 378312
rect 252374 378800 252430 378856
rect 253570 378528 253626 378584
rect 258354 378528 258410 378584
rect 260930 378528 260986 378584
rect 252374 378392 252430 378448
rect 250626 378256 250682 378312
rect 270958 380568 271014 380624
rect 268658 379380 268660 379400
rect 268660 379380 268712 379400
rect 268712 379380 268714 379400
rect 268658 379344 268714 379380
rect 263598 378528 263654 378584
rect 265898 378528 265954 378584
rect 268106 378528 268162 378584
rect 262862 378392 262918 378448
rect 262770 378256 262826 378312
rect 266358 378256 266414 378312
rect 267554 378256 267610 378312
rect 271050 379364 271106 379400
rect 271050 379344 271052 379364
rect 271052 379344 271104 379364
rect 271104 379344 271106 379364
rect 272062 379344 272118 379400
rect 273258 379344 273314 379400
rect 274178 379344 274234 379400
rect 275650 379344 275706 379400
rect 276018 379344 276074 379400
rect 276938 379344 276994 379400
rect 285954 379344 286010 379400
rect 287702 379344 287758 379400
rect 290922 379344 290978 379400
rect 292670 379344 292726 379400
rect 273442 378528 273498 378584
rect 274638 378156 274640 378176
rect 274640 378156 274692 378176
rect 274692 378156 274694 378176
rect 274638 378120 274694 378156
rect 277858 379208 277914 379264
rect 278042 379208 278098 379264
rect 279146 379208 279202 379264
rect 280710 379208 280766 379264
rect 283010 379208 283066 379264
rect 295890 379344 295946 379400
rect 298466 379344 298522 379400
rect 300858 379344 300914 379400
rect 433430 574504 433486 574560
rect 433522 560360 433578 560416
rect 433614 546352 433670 546408
rect 433522 522552 433578 522608
rect 429198 520104 429254 520160
rect 434902 628088 434958 628144
rect 456798 627680 456854 627736
rect 436282 623328 436338 623384
rect 436190 613808 436246 613864
rect 436098 609048 436154 609104
rect 436098 604288 436154 604344
rect 434902 585248 434958 585304
rect 434810 532208 434866 532264
rect 434718 519968 434774 520024
rect 397458 516704 397514 516760
rect 302790 379344 302846 379400
rect 305826 379344 305882 379400
rect 310978 379344 311034 379400
rect 313370 379364 313426 379400
rect 313370 379344 313372 379364
rect 313372 379344 313424 379364
rect 313424 379344 313426 379364
rect 315762 379380 315764 379400
rect 315764 379380 315816 379400
rect 315816 379380 315818 379400
rect 315762 379344 315818 379380
rect 317418 379344 317474 379400
rect 323306 379344 323362 379400
rect 325974 379344 326030 379400
rect 343454 379344 343510 379400
rect 320914 378528 320970 378584
rect 343178 378392 343234 378448
rect 338486 358828 338542 358864
rect 338486 358808 338488 358828
rect 338488 358808 338540 358828
rect 338540 358808 338542 358828
rect 339866 358808 339922 358864
rect 351734 358808 351790 358864
rect 273166 273808 273222 273864
rect 266358 273556 266414 273592
rect 266358 273536 266360 273556
rect 266360 273536 266412 273556
rect 266412 273536 266414 273556
rect 269762 273536 269818 273592
rect 271142 273536 271198 273592
rect 283470 273536 283526 273592
rect 273258 273400 273314 273456
rect 298466 273012 298522 273048
rect 298466 272992 298468 273012
rect 298468 272992 298520 273012
rect 298520 272992 298522 273012
rect 285954 272856 286010 272912
rect 288162 272856 288218 272912
rect 290922 272876 290978 272912
rect 290922 272856 290924 272876
rect 290924 272856 290976 272876
rect 290976 272856 290978 272876
rect 293314 272856 293370 272912
rect 295890 272892 295892 272912
rect 295892 272892 295944 272912
rect 295944 272892 295946 272912
rect 295890 272856 295946 272892
rect 300858 272740 300914 272776
rect 300858 272720 300860 272740
rect 300860 272720 300912 272740
rect 300912 272720 300914 272740
rect 303434 272720 303490 272776
rect 310978 272604 311034 272640
rect 310978 272584 310980 272604
rect 310980 272584 311032 272604
rect 311032 272584 311034 272604
rect 320914 272584 320970 272640
rect 265162 272176 265218 272232
rect 263598 271768 263654 271824
rect 260838 271380 260894 271416
rect 260838 271360 260840 271380
rect 260840 271360 260892 271380
rect 260892 271360 260894 271380
rect 258262 271224 258318 271280
rect 264978 271244 265034 271280
rect 264978 271224 264980 271244
rect 264980 271224 265032 271244
rect 265032 271224 265034 271244
rect 247038 271088 247094 271144
rect 252558 271088 252614 271144
rect 255318 271108 255374 271144
rect 255318 271088 255320 271108
rect 255320 271088 255372 271108
rect 255372 271088 255374 271108
rect 253938 270816 253994 270872
rect 244370 270680 244426 270736
rect 251270 270680 251326 270736
rect 235998 270544 236054 270600
rect 237378 270544 237434 270600
rect 242898 270544 242954 270600
rect 244278 270544 244334 270600
rect 245658 270544 245714 270600
rect 247038 270544 247094 270600
rect 248510 270544 248566 270600
rect 249798 270544 249854 270600
rect 251178 270544 251234 270600
rect 252558 270544 252614 270600
rect 255318 270680 255374 270736
rect 259550 270680 259606 270736
rect 256698 270544 256754 270600
rect 258078 270544 258134 270600
rect 259458 270544 259514 270600
rect 260838 270544 260894 270600
rect 262218 270544 262274 270600
rect 263598 270544 263654 270600
rect 270498 271768 270554 271824
rect 271878 271768 271934 271824
rect 276018 271768 276074 271824
rect 277950 271768 278006 271824
rect 280158 271768 280214 271824
rect 307758 271788 307814 271824
rect 307758 271768 307760 271788
rect 307760 271768 307812 271788
rect 307812 271768 307814 271788
rect 267830 271360 267886 271416
rect 266358 270544 266414 270600
rect 268198 270544 268254 270600
rect 276018 271532 276020 271552
rect 276020 271532 276072 271552
rect 276072 271532 276074 271552
rect 276018 271496 276074 271532
rect 343546 271804 343548 271824
rect 343548 271804 343600 271824
rect 343600 271804 343602 271824
rect 343546 271768 343602 271804
rect 343546 271360 343602 271416
rect 275926 271224 275982 271280
rect 278686 271244 278742 271280
rect 278686 271224 278688 271244
rect 278688 271224 278740 271244
rect 278740 271224 278742 271244
rect 313278 271088 313334 271144
rect 280066 270816 280122 270872
rect 340786 253408 340842 253464
rect 351826 253172 351828 253192
rect 351828 253172 351880 253192
rect 351880 253172 351882 253192
rect 351826 253136 351882 253172
rect 339406 253000 339462 253056
rect 288070 166640 288126 166696
rect 288254 166640 288310 166696
rect 291014 166640 291070 166696
rect 260930 166368 260986 166424
rect 265898 166368 265954 166424
rect 288070 166368 288126 166424
rect 293314 166388 293370 166424
rect 293314 166368 293316 166388
rect 293316 166368 293368 166388
rect 293368 166368 293370 166388
rect 298466 166368 298522 166424
rect 285954 166232 286010 166288
rect 236090 165552 236146 165608
rect 238758 165552 238814 165608
rect 242898 165552 242954 165608
rect 247130 165552 247186 165608
rect 255318 165552 255374 165608
rect 258170 165552 258226 165608
rect 260838 165552 260894 165608
rect 277398 165552 277454 165608
rect 280158 165552 280214 165608
rect 283378 165552 283434 165608
rect 300858 165552 300914 165608
rect 308218 165552 308274 165608
rect 320914 165552 320970 165608
rect 325882 165572 325938 165608
rect 325882 165552 325884 165572
rect 325884 165552 325936 165572
rect 325936 165552 325938 165572
rect 235998 164192 236054 164248
rect 237378 164192 237434 164248
rect 220818 145832 220874 145888
rect 240138 164192 240194 164248
rect 241518 164192 241574 164248
rect 247038 164872 247094 164928
rect 244278 164328 244334 164384
rect 244370 164192 244426 164248
rect 245658 164192 245714 164248
rect 249798 164892 249854 164928
rect 249798 164872 249800 164892
rect 249800 164872 249852 164892
rect 249852 164872 249854 164892
rect 252558 164872 252614 164928
rect 258078 164872 258134 164928
rect 251270 164328 251326 164384
rect 248418 164192 248474 164248
rect 249890 164192 249946 164248
rect 251178 164192 251234 164248
rect 237378 145560 237434 145616
rect 252650 164192 252706 164248
rect 253938 164192 253994 164248
rect 255410 164192 255466 164248
rect 256698 164192 256754 164248
rect 259550 164328 259606 164384
rect 259458 164192 259514 164248
rect 264978 165144 265034 165200
rect 267738 165164 267794 165200
rect 267738 165144 267740 165164
rect 267740 165144 267792 165164
rect 267792 165144 267794 165164
rect 263506 164192 263562 164248
rect 263782 164192 263838 164248
rect 271878 165144 271934 165200
rect 274822 165144 274878 165200
rect 276018 165144 276074 165200
rect 280066 165144 280122 165200
rect 267646 164328 267702 164384
rect 266358 164192 266414 164248
rect 267738 164192 267794 164248
rect 263598 145968 263654 146024
rect 269118 164192 269174 164248
rect 270498 164192 270554 164248
rect 273442 165028 273498 165064
rect 273442 165008 273444 165028
rect 273444 165008 273496 165028
rect 273496 165008 273498 165028
rect 273810 164328 273866 164384
rect 274546 164192 274602 164248
rect 269118 146240 269174 146296
rect 277306 164192 277362 164248
rect 278042 164192 278098 164248
rect 278042 148960 278098 149016
rect 278686 148960 278742 149016
rect 278686 148280 278742 148336
rect 267830 146104 267886 146160
rect 267738 145832 267794 145888
rect 343270 165572 343326 165608
rect 343270 165552 343272 165572
rect 343272 165552 343324 165572
rect 343324 165552 343326 165572
rect 343454 165552 343510 165608
rect 308218 163920 308274 163976
rect 338486 144880 338542 144936
rect 340234 144880 340290 144936
rect 351642 144880 351698 144936
rect 235998 59744 236054 59800
rect 237102 59744 237158 59800
rect 255870 59744 255926 59800
rect 256974 59744 257030 59800
rect 262862 59744 262918 59800
rect 260654 59608 260710 59664
rect 259458 59336 259514 59392
rect 308494 59608 308550 59664
rect 315854 59608 315910 59664
rect 261666 59336 261722 59392
rect 279238 59200 279294 59256
rect 290922 59200 290978 59256
rect 300858 59200 300914 59256
rect 320914 59200 320970 59256
rect 325882 59200 325938 59256
rect 237378 57840 237434 57896
rect 239218 57840 239274 57896
rect 240138 57840 240194 57896
rect 241610 57840 241666 57896
rect 242898 57840 242954 57896
rect 244370 57840 244426 57896
rect 245290 57840 245346 57896
rect 245658 57840 245714 57896
rect 247682 57840 247738 57896
rect 248418 57840 248474 57896
rect 250074 57840 250130 57896
rect 250994 57840 251050 57896
rect 264978 57840 265034 57896
rect 271050 57840 271106 57896
rect 271878 57840 271934 57896
rect 273258 57840 273314 57896
rect 274638 57840 274694 57896
rect 276938 57840 276994 57896
rect 287610 57840 287666 57896
rect 293314 57840 293370 57896
rect 295890 57840 295946 57896
rect 298098 57840 298154 57896
rect 303434 57840 303490 57896
rect 305826 57840 305882 57896
rect 310978 57840 311034 57896
rect 313370 57860 313426 57896
rect 313370 57840 313372 57860
rect 313372 57840 313424 57860
rect 313424 57840 313426 57860
rect 258354 57704 258410 57760
rect 263598 57704 263654 57760
rect 250994 57432 251050 57488
rect 251178 57432 251234 57488
rect 251914 57432 251970 57488
rect 252558 57432 252614 57488
rect 253938 57432 253994 57488
rect 266450 57704 266506 57760
rect 268474 57704 268530 57760
rect 269118 57704 269174 57760
rect 266358 57432 266414 57488
rect 273350 57704 273406 57760
rect 269118 54984 269174 55040
rect 318246 57840 318302 57896
rect 323306 57876 323308 57896
rect 323308 57876 323360 57896
rect 323360 57876 323362 57896
rect 323306 57840 323362 57876
rect 343178 57876 343180 57896
rect 343180 57876 343232 57896
rect 343232 57876 343234 57896
rect 343178 57840 343234 57876
rect 343454 57860 343510 57896
rect 357438 148960 357494 149016
rect 358818 460128 358874 460184
rect 358910 400288 358966 400344
rect 359002 398112 359058 398168
rect 359094 394032 359150 394088
rect 358910 353096 358966 353152
rect 358818 291760 358874 291816
rect 359278 292712 359334 292768
rect 359186 290944 359242 291000
rect 359094 287544 359150 287600
rect 358910 246200 358966 246256
rect 358818 184864 358874 184920
rect 359830 396752 359886 396808
rect 359922 395256 359978 395312
rect 359738 371864 359794 371920
rect 359922 371864 359978 371920
rect 359554 292712 359610 292768
rect 359462 291760 359518 291816
rect 359738 288768 359794 288824
rect 359278 186360 359334 186416
rect 359462 186360 359518 186416
rect 359370 184864 359426 184920
rect 359186 183368 359242 183424
rect 359094 182008 359150 182064
rect 359002 180648 359058 180704
rect 359002 179424 359058 179480
rect 358910 139304 358966 139360
rect 359278 179424 359334 179480
rect 359186 76880 359242 76936
rect 359094 75384 359150 75440
rect 359554 182008 359610 182064
rect 359462 79872 359518 79928
rect 359370 78240 359426 78296
rect 359278 74024 359334 74080
rect 343454 57840 343456 57860
rect 343456 57840 343508 57860
rect 343508 57840 343510 57860
rect 365626 379480 365682 379536
rect 365534 379072 365590 379128
rect 366362 472640 366418 472696
rect 274638 55120 274694 55176
rect 136454 3984 136510 4040
rect 132958 3440 133014 3496
rect 129370 3304 129426 3360
rect 140042 3848 140098 3904
rect 147126 3712 147182 3768
rect 143538 3168 143594 3224
rect 150622 3576 150678 3632
rect 369766 273400 369822 273456
rect 369306 164600 369362 164656
rect 370318 145696 370374 145752
rect 369766 145560 369822 145616
rect 371146 379208 371202 379264
rect 371146 378664 371202 378720
rect 371146 376760 371202 376816
rect 371606 378120 371662 378176
rect 371698 269864 371754 269920
rect 373170 378936 373226 378992
rect 373170 378664 373226 378720
rect 372986 269184 373042 269240
rect 372250 146104 372306 146160
rect 374274 381520 374330 381576
rect 373538 270952 373594 271008
rect 373538 269184 373594 269240
rect 374366 271224 374422 271280
rect 375194 381520 375250 381576
rect 375010 378800 375066 378856
rect 376022 165280 376078 165336
rect 376390 380840 376446 380896
rect 376298 271496 376354 271552
rect 376942 417832 376998 417888
rect 377034 411984 377090 412040
rect 377034 410896 377090 410952
rect 376942 390904 376998 390960
rect 376942 389272 376998 389328
rect 376942 389000 376998 389056
rect 376482 270272 376538 270328
rect 376666 375128 376722 375184
rect 377770 416880 377826 416936
rect 377678 414724 377734 414760
rect 377678 414704 377680 414724
rect 377680 414704 377732 414724
rect 377732 414704 377734 414724
rect 377586 411984 377642 412040
rect 377402 409148 377458 409184
rect 377402 409128 377404 409148
rect 377404 409128 377456 409148
rect 377456 409128 377458 409148
rect 376942 310936 376998 310992
rect 376758 282104 376814 282160
rect 376942 284008 376998 284064
rect 376942 282240 376998 282296
rect 377126 302096 377182 302152
rect 377034 204176 377090 204232
rect 376942 203904 376998 203960
rect 377034 202952 377090 203008
rect 376942 201320 376998 201376
rect 376942 176976 376998 177032
rect 376942 175344 376998 175400
rect 376942 175072 376998 175128
rect 377310 309984 377366 310040
rect 377770 413752 377826 413808
rect 377678 307808 377734 307864
rect 377586 304952 377642 305008
rect 377494 303864 377550 303920
rect 377402 252492 377404 252512
rect 377404 252492 377456 252512
rect 377456 252492 377458 252512
rect 377402 252456 377458 252492
rect 377310 204176 377366 204232
rect 377310 203904 377366 203960
rect 377218 198736 377274 198792
rect 377126 195200 377182 195256
rect 377034 95920 377090 95976
rect 376942 93744 376998 93800
rect 378046 409128 378102 409184
rect 377954 374720 378010 374776
rect 377862 309984 377918 310040
rect 377770 306720 377826 306776
rect 377770 304952 377826 305008
rect 377678 201320 377734 201376
rect 377678 200776 377734 200832
rect 378046 302096 378102 302152
rect 377862 199824 377918 199880
rect 377862 198736 377918 198792
rect 377678 198056 377734 198112
rect 377586 196968 377642 197024
rect 377494 145560 377550 145616
rect 377310 96872 377366 96928
rect 377218 92792 377274 92848
rect 376942 69944 376998 70000
rect 376942 68332 376998 68368
rect 376942 68312 376944 68332
rect 376944 68312 376996 68332
rect 376996 68312 376998 68332
rect 377862 196968 377918 197024
rect 377770 195200 377826 195256
rect 377678 91024 377734 91080
rect 378414 146240 378470 146296
rect 378690 270408 378746 270464
rect 436834 599528 436890 599584
rect 436282 580488 436338 580544
rect 436190 536968 436246 537024
rect 436374 570288 436430 570344
rect 436466 565528 436522 565584
rect 436282 527448 436338 527504
rect 436558 556008 436614 556064
rect 436650 551248 436706 551304
rect 436742 541728 436798 541784
rect 580170 683848 580226 683904
rect 477130 627816 477186 627872
rect 488722 627816 488778 627872
rect 506754 627816 506810 627872
rect 457718 621560 457774 621616
rect 457626 615440 457682 615496
rect 580170 630808 580226 630864
rect 512182 624960 512238 625016
rect 512090 618840 512146 618896
rect 511998 612040 512054 612096
rect 457534 609320 457590 609376
rect 511998 605920 512054 605976
rect 457626 602520 457682 602576
rect 457534 596400 457590 596456
rect 457442 590280 457498 590336
rect 457442 584160 457498 584216
rect 436374 522416 436430 522472
rect 378782 165416 378838 165472
rect 379058 271632 379114 271688
rect 506478 515344 506534 515400
rect 483018 490456 483074 490512
rect 512182 599800 512238 599856
rect 512090 593680 512146 593736
rect 511998 487736 512054 487792
rect 512274 587560 512330 587616
rect 513010 580760 513066 580816
rect 580262 577632 580318 577688
rect 512090 479440 512146 479496
rect 457534 478080 457590 478136
rect 498474 466556 498476 466576
rect 498476 466556 498528 466576
rect 498528 466556 498530 466576
rect 498474 466520 498530 466556
rect 499762 466540 499818 466576
rect 499762 466520 499764 466540
rect 499764 466520 499816 466540
rect 499816 466520 499818 466540
rect 510894 466540 510950 466576
rect 510894 466520 510896 466540
rect 510896 466520 510948 466540
rect 510948 466520 510950 466540
rect 379610 382336 379666 382392
rect 421102 380704 421158 380760
rect 422850 380704 422906 380760
rect 430946 380704 431002 380760
rect 433614 380704 433670 380760
rect 436006 380704 436062 380760
rect 438490 380704 438546 380760
rect 440882 380704 440938 380760
rect 443458 380704 443514 380760
rect 408682 380568 408738 380624
rect 413466 380568 413522 380624
rect 419446 380568 419502 380624
rect 434350 380568 434406 380624
rect 379610 375264 379666 375320
rect 379426 273400 379482 273456
rect 379242 269864 379298 269920
rect 379242 269320 379298 269376
rect 379058 264968 379114 265024
rect 378414 145968 378470 146024
rect 377954 145832 378010 145888
rect 377954 145560 378010 145616
rect 377862 89936 377918 89992
rect 377770 88168 377826 88224
rect 379794 271088 379850 271144
rect 379702 270408 379758 270464
rect 379702 269728 379758 269784
rect 445942 380568 445998 380624
rect 396078 379344 396134 379400
rect 397090 379344 397146 379400
rect 403622 379344 403678 379400
rect 405830 379344 405886 379400
rect 407578 379344 407634 379400
rect 408314 379364 408370 379400
rect 408314 379344 408316 379364
rect 408316 379344 408368 379364
rect 408368 379344 408370 379364
rect 402978 379208 403034 379264
rect 405370 379208 405426 379264
rect 411258 379344 411314 379400
rect 412362 379344 412418 379400
rect 413098 379344 413154 379400
rect 414570 379344 414626 379400
rect 423402 379344 423458 379400
rect 426438 379344 426494 379400
rect 426622 379344 426678 379400
rect 435730 379380 435732 379400
rect 435732 379380 435784 379400
rect 435784 379380 435786 379400
rect 435730 379344 435786 379380
rect 439042 379344 439098 379400
rect 447506 379344 447562 379400
rect 451002 379344 451058 379400
rect 452750 379344 452806 379400
rect 455602 379344 455658 379400
rect 458362 379344 458418 379400
rect 460938 379344 460994 379400
rect 463514 379344 463570 379400
rect 474830 379344 474886 379400
rect 410062 379208 410118 379264
rect 409970 378120 410026 378176
rect 415766 379208 415822 379264
rect 416042 379208 416098 379264
rect 418250 378664 418306 378720
rect 416962 378528 417018 378584
rect 418158 378120 418214 378176
rect 419630 378120 419686 378176
rect 421746 378120 421802 378176
rect 425978 378664 426034 378720
rect 423954 378120 424010 378176
rect 425150 378120 425206 378176
rect 437754 379208 437810 379264
rect 427910 378664 427966 378720
rect 436466 378528 436522 378584
rect 431130 378256 431186 378312
rect 428278 378120 428334 378176
rect 429290 378120 429346 378176
rect 432234 378120 432290 378176
rect 473450 379208 473506 379264
rect 465078 379072 465134 379128
rect 463514 377984 463570 378040
rect 467930 378800 467986 378856
rect 470874 378800 470930 378856
rect 480534 379208 480590 379264
rect 503074 379208 503130 379264
rect 503534 379208 503590 379264
rect 477590 378936 477646 378992
rect 483386 378936 483442 378992
rect 483386 376624 483442 376680
rect 498934 358808 498990 358864
rect 500774 358808 500830 358864
rect 510894 358828 510950 358864
rect 510894 358808 510896 358828
rect 510896 358808 510948 358828
rect 510948 358808 510950 358828
rect 421102 273536 421158 273592
rect 422850 273536 422906 273592
rect 427634 273536 427690 273592
rect 445942 273536 445998 273592
rect 423402 272992 423458 273048
rect 425242 272992 425298 273048
rect 425978 273028 425980 273048
rect 425980 273028 426032 273048
rect 426032 273028 426034 273048
rect 425978 272992 426034 273028
rect 428186 273012 428242 273048
rect 428186 272992 428188 273012
rect 428188 272992 428240 273012
rect 428240 272992 428242 273012
rect 468482 272992 468538 273048
rect 470874 272856 470930 272912
rect 478418 272876 478474 272912
rect 478418 272856 478420 272876
rect 478420 272856 478472 272876
rect 478472 272856 478474 272876
rect 473450 272740 473506 272776
rect 473450 272720 473452 272740
rect 473452 272720 473504 272740
rect 473504 272720 473506 272740
rect 480810 272720 480866 272776
rect 475842 272604 475898 272640
rect 475842 272584 475844 272604
rect 475844 272584 475896 272604
rect 475896 272584 475898 272604
rect 485962 272584 486018 272640
rect 401690 272176 401746 272232
rect 415858 272176 415914 272232
rect 416042 272176 416098 272232
rect 455786 272176 455842 272232
rect 390558 269320 390614 269376
rect 388442 269184 388498 269240
rect 397458 270544 397514 270600
rect 398838 270544 398894 270600
rect 400218 270544 400274 270600
rect 409878 271088 409934 271144
rect 412730 271088 412786 271144
rect 418158 271108 418214 271144
rect 418158 271088 418160 271108
rect 418160 271088 418212 271108
rect 418212 271088 418214 271108
rect 405738 270816 405794 270872
rect 402978 270544 403034 270600
rect 403622 270544 403678 270600
rect 404358 270544 404414 270600
rect 411350 270680 411406 270736
rect 407118 270544 407174 270600
rect 408498 270544 408554 270600
rect 409878 270544 409934 270600
rect 411258 270544 411314 270600
rect 413006 270544 413062 270600
rect 414018 270544 414074 270600
rect 416778 270544 416834 270600
rect 418158 270544 418214 270600
rect 419538 270544 419594 270600
rect 420918 270544 420974 270600
rect 427818 271768 427874 271824
rect 430578 271768 430634 271824
rect 432050 271768 432106 271824
rect 433338 271768 433394 271824
rect 434718 271768 434774 271824
rect 437478 271768 437534 271824
rect 442998 271768 443054 271824
rect 447138 271768 447194 271824
rect 449898 271768 449954 271824
rect 452658 271768 452714 271824
rect 458178 271804 458180 271824
rect 458180 271804 458232 271824
rect 458232 271804 458234 271824
rect 433338 271360 433394 271416
rect 458178 271768 458234 271804
rect 503626 271632 503682 271688
rect 440238 271360 440294 271416
rect 440146 271224 440202 271280
rect 503626 271244 503682 271280
rect 503626 271224 503628 271244
rect 503628 271224 503680 271244
rect 503680 271224 503682 271244
rect 434718 270816 434774 270872
rect 436098 270816 436154 270872
rect 437478 270816 437534 270872
rect 429198 270680 429254 270736
rect 434810 270680 434866 270736
rect 500866 253308 500868 253328
rect 500868 253308 500920 253328
rect 500920 253308 500922 253328
rect 500866 253272 500922 253308
rect 499210 252728 499266 252784
rect 510894 252612 510950 252648
rect 510894 252592 510896 252612
rect 510896 252592 510948 252612
rect 510948 252592 510950 252612
rect 418434 166812 418436 166832
rect 418436 166812 418488 166832
rect 418488 166812 418490 166832
rect 418434 166776 418490 166812
rect 421010 166796 421066 166832
rect 421010 166776 421012 166796
rect 421012 166776 421064 166796
rect 421064 166776 421066 166796
rect 428278 166776 428334 166832
rect 430946 166776 431002 166832
rect 433614 166776 433670 166832
rect 473450 166776 473506 166832
rect 475842 166776 475898 166832
rect 478418 166776 478474 166832
rect 480902 166776 480958 166832
rect 434350 166504 434406 166560
rect 423402 166252 423458 166288
rect 423402 166232 423404 166252
rect 423404 166232 423456 166252
rect 423456 166232 423458 166252
rect 483386 166640 483442 166696
rect 485962 166640 486018 166696
rect 503258 166504 503314 166560
rect 397458 165552 397514 165608
rect 401598 165552 401654 165608
rect 404358 165552 404414 165608
rect 407118 165552 407174 165608
rect 415490 165552 415546 165608
rect 416042 165552 416098 165608
rect 418710 165552 418766 165608
rect 423678 165552 423734 165608
rect 426530 165552 426586 165608
rect 429658 165552 429714 165608
rect 435086 165552 435142 165608
rect 435914 165552 435970 165608
rect 437938 165552 437994 165608
rect 438490 165552 438546 165608
rect 440146 165552 440202 165608
rect 440882 165552 440938 165608
rect 443458 165552 443514 165608
rect 445850 165552 445906 165608
rect 447322 165552 447378 165608
rect 449898 165552 449954 165608
rect 452658 165552 452714 165608
rect 455418 165552 455474 165608
rect 458362 165572 458418 165608
rect 458362 165552 458364 165572
rect 458364 165552 458416 165572
rect 458416 165552 458418 165572
rect 396170 164328 396226 164384
rect 396078 164192 396134 164248
rect 398838 164192 398894 164248
rect 400218 164192 400274 164248
rect 403070 164328 403126 164384
rect 402978 164192 403034 164248
rect 412638 164892 412694 164928
rect 412638 164872 412640 164892
rect 412640 164872 412692 164892
rect 412692 164872 412694 164892
rect 409878 164756 409934 164792
rect 409878 164736 409880 164756
rect 409880 164736 409932 164756
rect 409932 164736 409934 164756
rect 411350 164328 411406 164384
rect 405738 164192 405794 164248
rect 407210 164192 407266 164248
rect 408498 164192 408554 164248
rect 409970 164192 410026 164248
rect 411258 164192 411314 164248
rect 412638 164192 412694 164248
rect 414018 164192 414074 164248
rect 416778 164192 416834 164248
rect 418158 164192 418214 164248
rect 420918 164464 420974 164520
rect 419538 164192 419594 164248
rect 422298 164192 422354 164248
rect 415490 145968 415546 146024
rect 425058 164192 425114 164248
rect 426438 164192 426494 164248
rect 423678 145832 423734 145888
rect 429106 164192 429162 164248
rect 432234 165008 432290 165064
rect 430578 164464 430634 164520
rect 425058 145696 425114 145752
rect 436190 164872 436246 164928
rect 434626 164192 434682 164248
rect 503350 165552 503406 165608
rect 518898 459584 518954 459640
rect 519450 459584 519506 459640
rect 519082 400288 519138 400344
rect 518990 398112 519046 398168
rect 440238 148280 440294 148336
rect 429198 145560 429254 145616
rect 510618 145424 510674 145480
rect 498658 144880 498714 144936
rect 500222 144880 500278 144936
rect 396078 59744 396134 59800
rect 397090 59764 397146 59800
rect 397090 59744 397092 59764
rect 397092 59744 397144 59764
rect 397144 59744 397146 59764
rect 403070 59744 403126 59800
rect 416962 59744 417018 59800
rect 422850 59744 422906 59800
rect 423954 59744 424010 59800
rect 404174 59608 404230 59664
rect 412546 59608 412602 59664
rect 410706 59336 410762 59392
rect 397458 57840 397514 57896
rect 399482 57840 399538 57896
rect 400218 57840 400274 57896
rect 401690 57840 401746 57896
rect 404358 57840 404414 57896
rect 405830 57840 405886 57896
rect 407210 57840 407266 57896
rect 408314 57840 408370 57896
rect 408682 57840 408738 57896
rect 409878 57840 409934 57896
rect 411350 57840 411406 57896
rect 411258 56888 411314 56944
rect 423494 59608 423550 59664
rect 414570 59356 414626 59392
rect 414570 59336 414572 59356
rect 414572 59336 414624 59356
rect 414624 59336 414626 59356
rect 416042 59336 416098 59392
rect 418158 59336 418214 59392
rect 419354 59336 419410 59392
rect 420642 59336 420698 59392
rect 421746 59336 421802 59392
rect 428186 59336 428242 59392
rect 475842 58928 475898 58984
rect 468482 58812 468538 58848
rect 468482 58792 468484 58812
rect 468484 58792 468536 58812
rect 468536 58792 468538 58812
rect 519174 396752 519230 396808
rect 519358 395256 519414 395312
rect 519266 394032 519322 394088
rect 519082 352960 519138 353016
rect 518898 292440 518954 292496
rect 518990 290264 519046 290320
rect 518898 186360 518954 186416
rect 415490 57840 415546 57896
rect 425242 57840 425298 57896
rect 426438 57840 426494 57896
rect 428554 57840 428610 57896
rect 429198 57840 429254 57896
rect 430578 57840 430634 57896
rect 432234 57840 432290 57896
rect 433522 57840 433578 57896
rect 434626 57840 434682 57896
rect 435914 57840 435970 57896
rect 436374 57840 436430 57896
rect 438490 57840 438546 57896
rect 445850 57840 445906 57896
rect 460938 57840 460994 57896
rect 465906 57840 465962 57896
rect 470874 57860 470930 57896
rect 470874 57840 470876 57860
rect 470876 57840 470928 57860
rect 470928 57840 470930 57860
rect 412546 56888 412602 56944
rect 412638 56752 412694 56808
rect 425242 55936 425298 55992
rect 426530 57160 426586 57216
rect 428554 56072 428610 56128
rect 430946 57160 431002 57216
rect 433154 57432 433210 57488
rect 433430 57432 433486 57488
rect 433154 57160 433210 57216
rect 434718 57432 434774 57488
rect 478418 57840 478474 57896
rect 485962 57876 485964 57896
rect 485964 57876 486016 57896
rect 486016 57876 486018 57896
rect 485962 57840 486018 57876
rect 503258 57876 503260 57896
rect 503260 57876 503312 57896
rect 503312 57876 503314 57896
rect 503258 57840 503314 57876
rect 503534 57860 503590 57896
rect 519174 288496 519230 288552
rect 519082 246200 519138 246256
rect 518990 183368 519046 183424
rect 518990 181872 519046 181928
rect 518898 79872 518954 79928
rect 580170 511264 580226 511320
rect 580262 458088 580318 458144
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 519450 352960 519506 353016
rect 519358 293800 519414 293856
rect 519266 287544 519322 287600
rect 519174 181872 519230 181928
rect 519450 292440 519506 292496
rect 519358 186360 519414 186416
rect 519542 290264 519598 290320
rect 580354 351872 580410 351928
rect 580262 325216 580318 325272
rect 519634 288496 519690 288552
rect 520186 288496 520242 288552
rect 580354 272176 580410 272232
rect 580262 232328 580318 232384
rect 580354 192480 580410 192536
rect 519450 184728 519506 184784
rect 520186 184728 520242 184784
rect 519358 183368 519414 183424
rect 519266 180648 519322 180704
rect 519082 139304 519138 139360
rect 518990 75384 519046 75440
rect 520094 183368 520150 183424
rect 580262 152632 580318 152688
rect 520186 79872 520242 79928
rect 519450 78240 519506 78296
rect 519358 76744 519414 76800
rect 519174 74160 519230 74216
rect 503534 57840 503536 57860
rect 503536 57840 503588 57860
rect 503588 57840 503590 57860
rect 437478 57432 437534 57488
rect 580446 112784 580502 112840
rect 580354 72936 580410 72992
rect 580262 33088 580318 33144
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect 324773 634946 324839 634949
rect 423857 634946 423923 634949
rect 324773 634944 423923 634946
rect 324773 634888 324778 634944
rect 324834 634888 423862 634944
rect 423918 634888 423923 634944
rect 324773 634886 423923 634888
rect 324773 634883 324839 634886
rect 423857 634883 423923 634886
rect 54334 632572 54340 632636
rect 54404 632634 54410 632636
rect 333053 632634 333119 632637
rect 54404 632632 333119 632634
rect 54404 632576 333058 632632
rect 333114 632576 333119 632632
rect 54404 632574 333119 632576
rect 54404 632572 54410 632574
rect 333053 632571 333119 632574
rect 53046 632436 53052 632500
rect 53116 632498 53122 632500
rect 351085 632498 351151 632501
rect 53116 632496 351151 632498
rect 53116 632440 351090 632496
rect 351146 632440 351151 632496
rect 53116 632438 351151 632440
rect 53116 632436 53122 632438
rect 351085 632435 351151 632438
rect 321093 632226 321159 632229
rect 321093 632224 325036 632226
rect -960 632090 480 632180
rect 321093 632168 321098 632224
rect 321154 632168 325036 632224
rect 321093 632166 325036 632168
rect 321093 632163 321159 632166
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect 57605 628690 57671 628693
rect 146293 628690 146359 628693
rect 237373 628690 237439 628693
rect 57605 628688 60106 628690
rect 57605 628632 57610 628688
rect 57666 628632 60106 628688
rect 57605 628630 60106 628632
rect 57605 628627 57671 628630
rect 60046 628592 60106 628630
rect 146293 628688 150082 628690
rect 146293 628632 146298 628688
rect 146354 628632 150082 628688
rect 146293 628630 150082 628632
rect 146293 628627 146359 628630
rect 150022 628592 150082 628630
rect 237373 628688 240242 628690
rect 237373 628632 237378 628688
rect 237434 628632 240242 628688
rect 237373 628630 240242 628632
rect 237373 628627 237439 628630
rect 240182 628592 240242 628630
rect 300853 628146 300919 628149
rect 434897 628146 434963 628149
rect 300718 628144 300919 628146
rect 300718 628088 300858 628144
rect 300914 628088 300919 628144
rect 300718 628086 300919 628088
rect 433780 628144 434963 628146
rect 433780 628088 434902 628144
rect 434958 628088 434963 628144
rect 433780 628086 434963 628088
rect 122833 628010 122899 628013
rect 211245 628010 211311 628013
rect 120766 628008 122899 628010
rect 120766 627952 122838 628008
rect 122894 627952 122899 628008
rect 120766 627950 122899 627952
rect 120766 627912 120826 627950
rect 122833 627947 122899 627950
rect 210742 628008 211311 628010
rect 210742 627952 211250 628008
rect 211306 627952 211311 628008
rect 210742 627950 211311 627952
rect 210742 627912 210802 627950
rect 211245 627947 211311 627950
rect 300718 627912 300778 628086
rect 300853 628083 300919 628086
rect 434897 628083 434963 628086
rect 476062 627812 476068 627876
rect 476132 627874 476138 627876
rect 477125 627874 477191 627877
rect 476132 627872 477191 627874
rect 476132 627816 477130 627872
rect 477186 627816 477191 627872
rect 476132 627814 477191 627816
rect 476132 627812 476138 627814
rect 477125 627811 477191 627814
rect 488574 627812 488580 627876
rect 488644 627874 488650 627876
rect 488717 627874 488783 627877
rect 488644 627872 488783 627874
rect 488644 627816 488722 627872
rect 488778 627816 488783 627872
rect 488644 627814 488783 627816
rect 488644 627812 488650 627814
rect 488717 627811 488783 627814
rect 506606 627812 506612 627876
rect 506676 627874 506682 627876
rect 506749 627874 506815 627877
rect 506676 627872 506815 627874
rect 506676 627816 506754 627872
rect 506810 627816 506815 627872
rect 506676 627814 506815 627816
rect 506676 627812 506682 627814
rect 506749 627811 506815 627814
rect 456793 627738 456859 627741
rect 456793 627736 460092 627738
rect 456793 627680 456798 627736
rect 456854 627680 460092 627736
rect 456793 627678 460092 627680
rect 456793 627675 456859 627678
rect 321553 627466 321619 627469
rect 321553 627464 325036 627466
rect 321553 627408 321558 627464
rect 321614 627408 325036 627464
rect 321553 627406 325036 627408
rect 321553 627403 321619 627406
rect 59261 625834 59327 625837
rect 59494 625834 60076 625870
rect 59261 625832 60076 625834
rect 59261 625776 59266 625832
rect 59322 625810 60076 625832
rect 148685 625834 148751 625837
rect 149470 625834 150052 625870
rect 148685 625832 150052 625834
rect 59322 625776 59554 625810
rect 59261 625774 59554 625776
rect 148685 625776 148690 625832
rect 148746 625810 150052 625832
rect 238293 625834 238359 625837
rect 239446 625834 240120 625870
rect 238293 625832 240120 625834
rect 148746 625776 149530 625810
rect 148685 625774 149530 625776
rect 238293 625776 238298 625832
rect 238354 625810 240120 625832
rect 238354 625776 239506 625810
rect 238293 625774 239506 625776
rect 59261 625771 59327 625774
rect 148685 625771 148751 625774
rect 238293 625771 238359 625774
rect 300945 625426 301011 625429
rect 300718 625424 301011 625426
rect 300718 625368 300950 625424
rect 301006 625368 301011 625424
rect 300718 625366 301011 625368
rect 123017 625290 123083 625293
rect 212717 625290 212783 625293
rect 120766 625288 123083 625290
rect 120766 625232 123022 625288
rect 123078 625232 123083 625288
rect 120766 625230 123083 625232
rect 120766 625192 120826 625230
rect 123017 625227 123083 625230
rect 210742 625288 212783 625290
rect 210742 625232 212722 625288
rect 212778 625232 212783 625288
rect 210742 625230 212783 625232
rect 210742 625192 210802 625230
rect 212717 625227 212783 625230
rect 300718 625192 300778 625366
rect 300945 625363 301011 625366
rect 512177 625018 512243 625021
rect 509956 625016 512243 625018
rect 509956 624960 512182 625016
rect 512238 624960 512243 625016
rect 509956 624958 512243 624960
rect 512177 624955 512243 624958
rect 436277 623386 436343 623389
rect 433780 623384 436343 623386
rect 433780 623328 436282 623384
rect 436338 623328 436343 623384
rect 433780 623326 436343 623328
rect 436277 623323 436343 623326
rect 321553 622706 321619 622709
rect 321553 622704 325036 622706
rect 321553 622648 321558 622704
rect 321614 622648 325036 622704
rect 321553 622646 325036 622648
rect 321553 622643 321619 622646
rect 57421 622434 57487 622437
rect 59494 622434 60076 622470
rect 57421 622432 60076 622434
rect 57421 622376 57426 622432
rect 57482 622410 60076 622432
rect 147305 622434 147371 622437
rect 149470 622434 150052 622470
rect 147305 622432 150052 622434
rect 57482 622376 59554 622410
rect 57421 622374 59554 622376
rect 147305 622376 147310 622432
rect 147366 622410 150052 622432
rect 237373 622434 237439 622437
rect 239446 622434 240120 622470
rect 237373 622432 240120 622434
rect 147366 622376 149530 622410
rect 147305 622374 149530 622376
rect 237373 622376 237378 622432
rect 237434 622410 240120 622432
rect 237434 622376 239506 622410
rect 237373 622374 239506 622376
rect 57421 622371 57487 622374
rect 147305 622371 147371 622374
rect 237373 622371 237439 622374
rect 120766 621210 120826 621792
rect 121821 621210 121887 621213
rect 120766 621208 121887 621210
rect 120766 621152 121826 621208
rect 121882 621152 121887 621208
rect 120766 621150 121887 621152
rect 210742 621210 210802 621792
rect 213269 621210 213335 621213
rect 210742 621208 213335 621210
rect 210742 621152 213274 621208
rect 213330 621152 213335 621208
rect 210742 621150 213335 621152
rect 300718 621210 300778 621792
rect 457713 621618 457779 621621
rect 457713 621616 460092 621618
rect 457713 621560 457718 621616
rect 457774 621560 460092 621616
rect 457713 621558 460092 621560
rect 457713 621555 457779 621558
rect 302877 621210 302943 621213
rect 300718 621208 302943 621210
rect 300718 621152 302882 621208
rect 302938 621152 302943 621208
rect 300718 621150 302943 621152
rect 121821 621147 121887 621150
rect 213269 621147 213335 621150
rect 302877 621147 302943 621150
rect 57513 619714 57579 619717
rect 59494 619714 60076 619750
rect 57513 619712 60076 619714
rect 57513 619656 57518 619712
rect 57574 619690 60076 619712
rect 146293 619714 146359 619717
rect 149470 619714 150052 619750
rect 146293 619712 150052 619714
rect 57574 619656 59554 619690
rect 57513 619654 59554 619656
rect 146293 619656 146298 619712
rect 146354 619690 150052 619712
rect 237373 619714 237439 619717
rect 239446 619714 240120 619750
rect 237373 619712 240120 619714
rect 146354 619656 149530 619690
rect 146293 619654 149530 619656
rect 237373 619656 237378 619712
rect 237434 619690 240120 619712
rect 237434 619656 239506 619690
rect 237373 619654 239506 619656
rect 57513 619651 57579 619654
rect 146293 619651 146359 619654
rect 237373 619651 237439 619654
rect -960 619020 480 619260
rect 433333 619170 433399 619173
rect 433333 619168 433442 619170
rect 433333 619112 433338 619168
rect 433394 619112 433442 619168
rect 433333 619107 433442 619112
rect 120766 618490 120826 619072
rect 121678 618490 121684 618492
rect 120766 618430 121684 618490
rect 121678 618428 121684 618430
rect 121748 618428 121754 618492
rect 210742 618490 210802 619072
rect 211429 618490 211495 618493
rect 210742 618488 211495 618490
rect 210742 618432 211434 618488
rect 211490 618432 211495 618488
rect 210742 618430 211495 618432
rect 300718 618490 300778 619072
rect 433382 618596 433442 619107
rect 512085 618898 512151 618901
rect 509956 618896 512151 618898
rect 509956 618840 512090 618896
rect 512146 618840 512151 618896
rect 509956 618838 512151 618840
rect 512085 618835 512151 618838
rect 301129 618490 301195 618493
rect 300718 618488 301195 618490
rect 300718 618432 301134 618488
rect 301190 618432 301195 618488
rect 300718 618430 301195 618432
rect 211429 618427 211495 618430
rect 301129 618427 301195 618430
rect 321553 617946 321619 617949
rect 321553 617944 325036 617946
rect 321553 617888 321558 617944
rect 321614 617888 325036 617944
rect 321553 617886 325036 617888
rect 321553 617883 321619 617886
rect 583520 617388 584960 617628
rect 58985 616314 59051 616317
rect 59494 616314 60076 616350
rect 58985 616312 60076 616314
rect 58985 616256 58990 616312
rect 59046 616290 60076 616312
rect 146293 616314 146359 616317
rect 149470 616314 150052 616350
rect 146293 616312 150052 616314
rect 59046 616256 59554 616290
rect 58985 616254 59554 616256
rect 146293 616256 146298 616312
rect 146354 616290 150052 616312
rect 237373 616314 237439 616317
rect 239446 616314 240120 616350
rect 237373 616312 240120 616314
rect 146354 616256 149530 616290
rect 146293 616254 149530 616256
rect 237373 616256 237378 616312
rect 237434 616290 240120 616312
rect 237434 616256 239506 616290
rect 237373 616254 239506 616256
rect 58985 616251 59051 616254
rect 146293 616251 146359 616254
rect 237373 616251 237439 616254
rect 120766 615634 120826 615672
rect 121729 615634 121795 615637
rect 120766 615632 121795 615634
rect 120766 615576 121734 615632
rect 121790 615576 121795 615632
rect 120766 615574 121795 615576
rect 210742 615634 210802 615672
rect 211153 615634 211219 615637
rect 210742 615632 211219 615634
rect 210742 615576 211158 615632
rect 211214 615576 211219 615632
rect 210742 615574 211219 615576
rect 300718 615634 300778 615672
rect 301037 615634 301103 615637
rect 300718 615632 301103 615634
rect 300718 615576 301042 615632
rect 301098 615576 301103 615632
rect 300718 615574 301103 615576
rect 121729 615571 121795 615574
rect 211153 615571 211219 615574
rect 301037 615571 301103 615574
rect 457621 615498 457687 615501
rect 457621 615496 460092 615498
rect 457621 615440 457626 615496
rect 457682 615440 460092 615496
rect 457621 615438 460092 615440
rect 457621 615435 457687 615438
rect 436185 613866 436251 613869
rect 433780 613864 436251 613866
rect 433780 613808 436190 613864
rect 436246 613808 436251 613864
rect 433780 613806 436251 613808
rect 436185 613803 436251 613806
rect 59169 613594 59235 613597
rect 59494 613594 60076 613630
rect 59169 613592 60076 613594
rect 59169 613536 59174 613592
rect 59230 613570 60076 613592
rect 146845 613594 146911 613597
rect 149470 613594 150052 613630
rect 146845 613592 150052 613594
rect 59230 613536 59554 613570
rect 59169 613534 59554 613536
rect 146845 613536 146850 613592
rect 146906 613570 150052 613592
rect 237373 613594 237439 613597
rect 239446 613594 240120 613630
rect 237373 613592 240120 613594
rect 146906 613536 149530 613570
rect 146845 613534 149530 613536
rect 237373 613536 237378 613592
rect 237434 613570 240120 613592
rect 237434 613536 239506 613570
rect 237373 613534 239506 613536
rect 59169 613531 59235 613534
rect 146845 613531 146911 613534
rect 237373 613531 237439 613534
rect 321553 613186 321619 613189
rect 321553 613184 325036 613186
rect 321553 613128 321558 613184
rect 321614 613128 325036 613184
rect 321553 613126 325036 613128
rect 321553 613123 321619 613126
rect 120766 612778 120826 612952
rect 123109 612778 123175 612781
rect 120766 612776 123175 612778
rect 120766 612720 123114 612776
rect 123170 612720 123175 612776
rect 120766 612718 123175 612720
rect 210742 612778 210802 612952
rect 211337 612778 211403 612781
rect 210742 612776 211403 612778
rect 210742 612720 211342 612776
rect 211398 612720 211403 612776
rect 210742 612718 211403 612720
rect 300718 612778 300778 612952
rect 301221 612778 301287 612781
rect 300718 612776 301287 612778
rect 300718 612720 301226 612776
rect 301282 612720 301287 612776
rect 300718 612718 301287 612720
rect 123109 612715 123175 612718
rect 211337 612715 211403 612718
rect 301221 612715 301287 612718
rect 511993 612098 512059 612101
rect 509956 612096 512059 612098
rect 509956 612040 511998 612096
rect 512054 612040 512059 612096
rect 509956 612038 512059 612040
rect 511993 612035 512059 612038
rect 59077 610194 59143 610197
rect 59494 610194 60076 610230
rect 59077 610192 60076 610194
rect 59077 610136 59082 610192
rect 59138 610170 60076 610192
rect 148501 610194 148567 610197
rect 149470 610194 150052 610230
rect 148501 610192 150052 610194
rect 59138 610136 59554 610170
rect 59077 610134 59554 610136
rect 148501 610136 148506 610192
rect 148562 610170 150052 610192
rect 237373 610194 237439 610197
rect 239446 610194 240120 610230
rect 237373 610192 240120 610194
rect 148562 610136 149530 610170
rect 148501 610134 149530 610136
rect 237373 610136 237378 610192
rect 237434 610170 240120 610192
rect 237434 610136 239506 610170
rect 237373 610134 239506 610136
rect 59077 610131 59143 610134
rect 148501 610131 148567 610134
rect 237373 610131 237439 610134
rect 120766 608970 120826 609552
rect 121913 608970 121979 608973
rect 120766 608968 121979 608970
rect 120766 608912 121918 608968
rect 121974 608912 121979 608968
rect 120766 608910 121979 608912
rect 210742 608970 210802 609552
rect 212809 608970 212875 608973
rect 210742 608968 212875 608970
rect 210742 608912 212814 608968
rect 212870 608912 212875 608968
rect 210742 608910 212875 608912
rect 300718 608970 300778 609552
rect 457529 609378 457595 609381
rect 457529 609376 460092 609378
rect 457529 609320 457534 609376
rect 457590 609320 460092 609376
rect 457529 609318 460092 609320
rect 457529 609315 457595 609318
rect 436093 609106 436159 609109
rect 433780 609104 436159 609106
rect 433780 609048 436098 609104
rect 436154 609048 436159 609104
rect 433780 609046 436159 609048
rect 436093 609043 436159 609046
rect 302417 608970 302483 608973
rect 300718 608968 302483 608970
rect 300718 608912 302422 608968
rect 302478 608912 302483 608968
rect 300718 608910 302483 608912
rect 121913 608907 121979 608910
rect 212809 608907 212875 608910
rect 302417 608907 302483 608910
rect 321553 608426 321619 608429
rect 321553 608424 325036 608426
rect 321553 608368 321558 608424
rect 321614 608368 325036 608424
rect 321553 608366 325036 608368
rect 321553 608363 321619 608366
rect 57789 607610 57855 607613
rect 147581 607610 147647 607613
rect 238937 607610 239003 607613
rect 57789 607608 59554 607610
rect 57789 607552 57794 607608
rect 57850 607566 59554 607608
rect 147581 607608 149530 607610
rect 57850 607552 60076 607566
rect 57789 607550 60076 607552
rect 57789 607547 57855 607550
rect 59494 607506 60076 607550
rect 147581 607552 147586 607608
rect 147642 607566 149530 607608
rect 238937 607608 239506 607610
rect 147642 607552 150052 607566
rect 147581 607550 150052 607552
rect 147581 607547 147647 607550
rect 149470 607506 150052 607550
rect 238937 607552 238942 607608
rect 238998 607552 239506 607608
rect 238937 607550 239506 607552
rect 238937 607547 239003 607550
rect 239446 607542 239506 607550
rect 239446 607482 240032 607542
rect 120766 606389 120826 606832
rect 120766 606384 120875 606389
rect 120766 606328 120814 606384
rect 120870 606328 120875 606384
rect 120766 606326 120875 606328
rect 210742 606386 210802 606832
rect 211613 606386 211679 606389
rect 210742 606384 211679 606386
rect 210742 606328 211618 606384
rect 211674 606328 211679 606384
rect 210742 606326 211679 606328
rect 300718 606386 300778 606832
rect 302969 606386 303035 606389
rect 300718 606384 303035 606386
rect 300718 606328 302974 606384
rect 303030 606328 303035 606384
rect 300718 606326 303035 606328
rect 120809 606323 120875 606326
rect 211613 606323 211679 606326
rect 302969 606323 303035 606326
rect -960 605964 480 606204
rect 511993 605978 512059 605981
rect 509956 605976 512059 605978
rect 509956 605920 511998 605976
rect 512054 605920 512059 605976
rect 509956 605918 512059 605920
rect 511993 605915 512059 605918
rect 436093 604346 436159 604349
rect 433780 604344 436159 604346
rect 433780 604288 436098 604344
rect 436154 604288 436159 604344
rect 433780 604286 436159 604288
rect 436093 604283 436159 604286
rect 146201 604210 146267 604213
rect 238017 604210 238083 604213
rect 146201 604208 149530 604210
rect 146201 604152 146206 604208
rect 146262 604166 149530 604208
rect 238017 604208 239506 604210
rect 146262 604152 150052 604166
rect 146201 604150 150052 604152
rect 146201 604147 146267 604150
rect 57881 604074 57947 604077
rect 59494 604074 60076 604110
rect 149470 604106 150052 604150
rect 238017 604152 238022 604208
rect 238078 604152 239506 604208
rect 238017 604150 239506 604152
rect 238017 604147 238083 604150
rect 239446 604142 239506 604150
rect 239446 604082 240032 604142
rect 57881 604072 60076 604074
rect 57881 604016 57886 604072
rect 57942 604050 60076 604072
rect 583520 604060 584960 604300
rect 57942 604016 59554 604050
rect 57881 604014 59554 604016
rect 57881 604011 57947 604014
rect 321553 603666 321619 603669
rect 321553 603664 325036 603666
rect 321553 603608 321558 603664
rect 321614 603608 325036 603664
rect 321553 603606 325036 603608
rect 321553 603603 321619 603606
rect 120766 603122 120826 603432
rect 123293 603122 123359 603125
rect 120766 603120 123359 603122
rect 120766 603064 123298 603120
rect 123354 603064 123359 603120
rect 120766 603062 123359 603064
rect 210742 603122 210802 603432
rect 212901 603122 212967 603125
rect 210742 603120 212967 603122
rect 210742 603064 212906 603120
rect 212962 603064 212967 603120
rect 210742 603062 212967 603064
rect 300718 603122 300778 603432
rect 302509 603122 302575 603125
rect 300718 603120 302575 603122
rect 300718 603064 302514 603120
rect 302570 603064 302575 603120
rect 300718 603062 302575 603064
rect 123293 603059 123359 603062
rect 212901 603059 212967 603062
rect 302509 603059 302575 603062
rect 457621 602578 457687 602581
rect 457621 602576 460092 602578
rect 457621 602520 457626 602576
rect 457682 602520 460092 602576
rect 457621 602518 460092 602520
rect 457621 602515 457687 602518
rect 58893 601354 58959 601357
rect 59494 601354 60076 601390
rect 58893 601352 60076 601354
rect 58893 601296 58898 601352
rect 58954 601330 60076 601352
rect 148593 601354 148659 601357
rect 149470 601354 150052 601390
rect 148593 601352 150052 601354
rect 58954 601296 59554 601330
rect 58893 601294 59554 601296
rect 148593 601296 148598 601352
rect 148654 601330 150052 601352
rect 237373 601354 237439 601357
rect 239446 601354 240120 601390
rect 237373 601352 240120 601354
rect 148654 601296 149530 601330
rect 148593 601294 149530 601296
rect 237373 601296 237378 601352
rect 237434 601330 240120 601352
rect 237434 601296 239506 601330
rect 237373 601294 239506 601296
rect 58893 601291 58959 601294
rect 148593 601291 148659 601294
rect 237373 601291 237439 601294
rect 120766 600402 120826 600712
rect 123201 600402 123267 600405
rect 120766 600400 123267 600402
rect 120766 600344 123206 600400
rect 123262 600344 123267 600400
rect 120766 600342 123267 600344
rect 210742 600402 210802 600712
rect 211521 600402 211587 600405
rect 210742 600400 211587 600402
rect 210742 600344 211526 600400
rect 211582 600344 211587 600400
rect 210742 600342 211587 600344
rect 300718 600402 300778 600712
rect 301313 600402 301379 600405
rect 300718 600400 301379 600402
rect 300718 600344 301318 600400
rect 301374 600344 301379 600400
rect 300718 600342 301379 600344
rect 123201 600339 123267 600342
rect 211521 600339 211587 600342
rect 301313 600339 301379 600342
rect 512177 599858 512243 599861
rect 509956 599856 512243 599858
rect 509956 599800 512182 599856
rect 512238 599800 512243 599856
rect 509956 599798 512243 599800
rect 512177 599795 512243 599798
rect 436829 599586 436895 599589
rect 433780 599584 436895 599586
rect 433780 599528 436834 599584
rect 436890 599528 436895 599584
rect 433780 599526 436895 599528
rect 436829 599523 436895 599526
rect 321553 598906 321619 598909
rect 321553 598904 325036 598906
rect 321553 598848 321558 598904
rect 321614 598848 325036 598904
rect 321553 598846 325036 598848
rect 321553 598843 321619 598846
rect 57329 597954 57395 597957
rect 59494 597954 60076 597990
rect 57329 597952 60076 597954
rect 57329 597896 57334 597952
rect 57390 597930 60076 597952
rect 146293 597954 146359 597957
rect 149470 597954 150052 597990
rect 146293 597952 150052 597954
rect 57390 597896 59554 597930
rect 57329 597894 59554 597896
rect 146293 597896 146298 597952
rect 146354 597930 150052 597952
rect 237373 597954 237439 597957
rect 239446 597954 240120 597990
rect 237373 597952 240120 597954
rect 146354 597896 149530 597930
rect 146293 597894 149530 597896
rect 237373 597896 237378 597952
rect 237434 597930 240120 597952
rect 237434 597896 239506 597930
rect 237373 597894 239506 597896
rect 57329 597891 57395 597894
rect 146293 597891 146359 597894
rect 237373 597891 237439 597894
rect 120766 596730 120826 597312
rect 124121 596730 124187 596733
rect 120766 596728 124187 596730
rect 120766 596672 124126 596728
rect 124182 596672 124187 596728
rect 120766 596670 124187 596672
rect 210742 596730 210802 597312
rect 214097 596730 214163 596733
rect 210742 596728 214163 596730
rect 210742 596672 214102 596728
rect 214158 596672 214163 596728
rect 210742 596670 214163 596672
rect 300718 596730 300778 597312
rect 302693 596730 302759 596733
rect 300718 596728 302759 596730
rect 300718 596672 302698 596728
rect 302754 596672 302759 596728
rect 300718 596670 302759 596672
rect 124121 596667 124187 596670
rect 214097 596667 214163 596670
rect 302693 596667 302759 596670
rect 457529 596458 457595 596461
rect 457529 596456 460092 596458
rect 457529 596400 457534 596456
rect 457590 596400 460092 596456
rect 457529 596398 460092 596400
rect 457529 596395 457595 596398
rect 57789 595234 57855 595237
rect 59494 595234 60076 595270
rect 57789 595232 60076 595234
rect 57789 595176 57794 595232
rect 57850 595210 60076 595232
rect 147121 595234 147187 595237
rect 149470 595234 150052 595270
rect 147121 595232 150052 595234
rect 57850 595176 59554 595210
rect 57789 595174 59554 595176
rect 147121 595176 147126 595232
rect 147182 595210 150052 595232
rect 237373 595234 237439 595237
rect 239446 595234 240120 595270
rect 237373 595232 240120 595234
rect 147182 595176 149530 595210
rect 147121 595174 149530 595176
rect 237373 595176 237378 595232
rect 237434 595210 240120 595232
rect 237434 595176 239506 595210
rect 237373 595174 239506 595176
rect 57789 595171 57855 595174
rect 147121 595171 147187 595174
rect 237373 595171 237439 595174
rect 436134 594826 436140 594828
rect 433780 594766 436140 594826
rect 436134 594764 436140 594766
rect 436204 594764 436210 594828
rect 120766 594010 120826 594592
rect 122005 594010 122071 594013
rect 120766 594008 122071 594010
rect 120766 593952 122010 594008
rect 122066 593952 122071 594008
rect 120766 593950 122071 593952
rect 210742 594010 210802 594592
rect 211705 594010 211771 594013
rect 210742 594008 211771 594010
rect 210742 593952 211710 594008
rect 211766 593952 211771 594008
rect 210742 593950 211771 593952
rect 300718 594010 300778 594592
rect 324221 594146 324287 594149
rect 324221 594144 325036 594146
rect 324221 594088 324226 594144
rect 324282 594088 325036 594144
rect 324221 594086 325036 594088
rect 324221 594083 324287 594086
rect 301405 594010 301471 594013
rect 300718 594008 301471 594010
rect 300718 593952 301410 594008
rect 301466 593952 301471 594008
rect 300718 593950 301471 593952
rect 122005 593947 122071 593950
rect 211705 593947 211771 593950
rect 301405 593947 301471 593950
rect 512085 593738 512151 593741
rect 509956 593736 512151 593738
rect 509956 593680 512090 593736
rect 512146 593680 512151 593736
rect 509956 593678 512151 593680
rect 512085 593675 512151 593678
rect -960 592908 480 593148
rect 57237 591834 57303 591837
rect 59494 591834 60076 591870
rect 57237 591832 60076 591834
rect 57237 591776 57242 591832
rect 57298 591810 60076 591832
rect 148409 591834 148475 591837
rect 149470 591834 150052 591870
rect 148409 591832 150052 591834
rect 57298 591776 59554 591810
rect 57237 591774 59554 591776
rect 148409 591776 148414 591832
rect 148470 591810 150052 591832
rect 237373 591834 237439 591837
rect 239446 591834 240120 591870
rect 237373 591832 240120 591834
rect 148470 591776 149530 591810
rect 148409 591774 149530 591776
rect 237373 591776 237378 591832
rect 237434 591810 240120 591832
rect 237434 591776 239506 591810
rect 237373 591774 239506 591776
rect 57237 591771 57303 591774
rect 148409 591771 148475 591774
rect 237373 591771 237439 591774
rect 121085 591222 121151 591225
rect 120796 591220 121151 591222
rect 120796 591164 121090 591220
rect 121146 591164 121151 591220
rect 120796 591162 121151 591164
rect 121085 591159 121151 591162
rect 210742 590746 210802 591192
rect 213085 590746 213151 590749
rect 210742 590744 213151 590746
rect 210742 590688 213090 590744
rect 213146 590688 213151 590744
rect 210742 590686 213151 590688
rect 300718 590746 300778 591192
rect 583520 590868 584960 591108
rect 302601 590746 302667 590749
rect 300718 590744 302667 590746
rect 300718 590688 302606 590744
rect 302662 590688 302667 590744
rect 300718 590686 302667 590688
rect 213085 590683 213151 590686
rect 302601 590683 302667 590686
rect 457437 590338 457503 590341
rect 457437 590336 460092 590338
rect 457437 590280 457442 590336
rect 457498 590280 460092 590336
rect 457437 590278 460092 590280
rect 457437 590275 457503 590278
rect 433382 589525 433442 590036
rect 433333 589520 433442 589525
rect 433333 589464 433338 589520
rect 433394 589464 433442 589520
rect 433333 589462 433442 589464
rect 433333 589459 433399 589462
rect 321553 589386 321619 589389
rect 321553 589384 325036 589386
rect 321553 589328 321558 589384
rect 321614 589328 325036 589384
rect 321553 589326 325036 589328
rect 321553 589323 321619 589326
rect 57145 589114 57211 589117
rect 59494 589114 60076 589150
rect 57145 589112 60076 589114
rect 57145 589056 57150 589112
rect 57206 589090 60076 589112
rect 147213 589114 147279 589117
rect 149470 589114 150052 589150
rect 147213 589112 150052 589114
rect 57206 589056 59554 589090
rect 57145 589054 59554 589056
rect 147213 589056 147218 589112
rect 147274 589090 150052 589112
rect 237373 589114 237439 589117
rect 239446 589114 240120 589150
rect 237373 589112 240120 589114
rect 147274 589056 149530 589090
rect 147213 589054 149530 589056
rect 237373 589056 237378 589112
rect 237434 589090 240120 589112
rect 237434 589056 239506 589090
rect 237373 589054 239506 589056
rect 57145 589051 57211 589054
rect 147213 589051 147279 589054
rect 237373 589051 237439 589054
rect 120766 588026 120826 588472
rect 122097 588026 122163 588029
rect 120766 588024 122163 588026
rect 120766 587968 122102 588024
rect 122158 587968 122163 588024
rect 120766 587966 122163 587968
rect 210742 588026 210802 588472
rect 212993 588026 213059 588029
rect 210742 588024 213059 588026
rect 210742 587968 212998 588024
rect 213054 587968 213059 588024
rect 210742 587966 213059 587968
rect 300718 588026 300778 588472
rect 302233 588026 302299 588029
rect 300718 588024 302299 588026
rect 300718 587968 302238 588024
rect 302294 587968 302299 588024
rect 300718 587966 302299 587968
rect 122097 587963 122163 587966
rect 212993 587963 213059 587966
rect 302233 587963 302299 587966
rect 512269 587618 512335 587621
rect 509956 587616 512335 587618
rect 509956 587560 512274 587616
rect 512330 587560 512335 587616
rect 509956 587558 512335 587560
rect 512269 587555 512335 587558
rect 58801 585714 58867 585717
rect 59494 585714 60076 585750
rect 58801 585712 60076 585714
rect 58801 585656 58806 585712
rect 58862 585690 60076 585712
rect 146293 585714 146359 585717
rect 149470 585714 150052 585750
rect 146293 585712 150052 585714
rect 58862 585656 59554 585690
rect 58801 585654 59554 585656
rect 146293 585656 146298 585712
rect 146354 585690 150052 585712
rect 237373 585714 237439 585717
rect 239446 585714 240120 585750
rect 237373 585712 240120 585714
rect 146354 585656 149530 585690
rect 146293 585654 149530 585656
rect 237373 585656 237378 585712
rect 237434 585690 240120 585712
rect 237434 585656 239506 585690
rect 237373 585654 239506 585656
rect 58801 585651 58867 585654
rect 146293 585651 146359 585654
rect 237373 585651 237439 585654
rect 434897 585306 434963 585309
rect 433780 585304 434963 585306
rect 433780 585248 434902 585304
rect 434958 585248 434963 585304
rect 433780 585246 434963 585248
rect 434897 585243 434963 585246
rect 120766 584490 120826 585072
rect 123385 584490 123451 584493
rect 120766 584488 123451 584490
rect 120766 584432 123390 584488
rect 123446 584432 123451 584488
rect 120766 584430 123451 584432
rect 210742 584490 210802 585072
rect 211797 584490 211863 584493
rect 210742 584488 211863 584490
rect 210742 584432 211802 584488
rect 211858 584432 211863 584488
rect 210742 584430 211863 584432
rect 300718 584490 300778 585072
rect 321553 584626 321619 584629
rect 321553 584624 325036 584626
rect 321553 584568 321558 584624
rect 321614 584568 325036 584624
rect 321553 584566 325036 584568
rect 321553 584563 321619 584566
rect 302785 584490 302851 584493
rect 300718 584488 302851 584490
rect 300718 584432 302790 584488
rect 302846 584432 302851 584488
rect 300718 584430 302851 584432
rect 123385 584427 123451 584430
rect 211797 584427 211863 584430
rect 302785 584427 302851 584430
rect 457437 584218 457503 584221
rect 457437 584216 460092 584218
rect 457437 584160 457442 584216
rect 457498 584160 460092 584216
rect 457437 584158 460092 584160
rect 457437 584155 457503 584158
rect 57053 582994 57119 582997
rect 59494 582994 60076 583030
rect 57053 582992 60076 582994
rect 57053 582936 57058 582992
rect 57114 582970 60076 582992
rect 146293 582994 146359 582997
rect 149470 582994 150052 583030
rect 146293 582992 150052 582994
rect 57114 582936 59554 582970
rect 57053 582934 59554 582936
rect 146293 582936 146298 582992
rect 146354 582970 150052 582992
rect 236729 582994 236795 582997
rect 239446 582994 240120 583030
rect 236729 582992 240120 582994
rect 146354 582936 149530 582970
rect 146293 582934 149530 582936
rect 236729 582936 236734 582992
rect 236790 582970 240120 582992
rect 236790 582936 239506 582970
rect 236729 582934 239506 582936
rect 57053 582931 57119 582934
rect 146293 582931 146359 582934
rect 236729 582931 236795 582934
rect 120766 581770 120826 582352
rect 123477 581770 123543 581773
rect 120766 581768 123543 581770
rect 120766 581712 123482 581768
rect 123538 581712 123543 581768
rect 120766 581710 123543 581712
rect 210742 581770 210802 582352
rect 212533 581770 212599 581773
rect 210742 581768 212599 581770
rect 210742 581712 212538 581768
rect 212594 581712 212599 581768
rect 210742 581710 212599 581712
rect 300718 581770 300778 582352
rect 301497 581770 301563 581773
rect 300718 581768 301563 581770
rect 300718 581712 301502 581768
rect 301558 581712 301563 581768
rect 300718 581710 301563 581712
rect 123477 581707 123543 581710
rect 212533 581707 212599 581710
rect 301497 581707 301563 581710
rect 513005 580818 513071 580821
rect 509956 580816 513071 580818
rect 509956 580760 513010 580816
rect 513066 580760 513071 580816
rect 509956 580758 513071 580760
rect 513005 580755 513071 580758
rect 436277 580546 436343 580549
rect 433780 580544 436343 580546
rect 433780 580488 436282 580544
rect 436338 580488 436343 580544
rect 433780 580486 436343 580488
rect 436277 580483 436343 580486
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 321553 579866 321619 579869
rect 321553 579864 325036 579866
rect 321553 579808 321558 579864
rect 321614 579808 325036 579864
rect 321553 579806 325036 579808
rect 321553 579803 321619 579806
rect 57421 579730 57487 579733
rect 146293 579730 146359 579733
rect 237373 579730 237439 579733
rect 57421 579728 59554 579730
rect 57421 579672 57426 579728
rect 57482 579686 59554 579728
rect 146293 579728 149530 579730
rect 57482 579672 60076 579686
rect 57421 579670 60076 579672
rect 57421 579667 57487 579670
rect 59494 579626 60076 579670
rect 146293 579672 146298 579728
rect 146354 579686 149530 579728
rect 237373 579728 239506 579730
rect 146354 579672 150052 579686
rect 146293 579670 150052 579672
rect 146293 579667 146359 579670
rect 149470 579626 150052 579670
rect 237373 579672 237378 579728
rect 237434 579672 239506 579728
rect 237373 579670 239506 579672
rect 237373 579667 237439 579670
rect 239446 579662 239506 579670
rect 239446 579602 240032 579662
rect 121177 578982 121243 578985
rect 120796 578980 121243 578982
rect 120796 578924 121182 578980
rect 121238 578924 121243 578980
rect 120796 578922 121243 578924
rect 121177 578919 121243 578922
rect 210742 578370 210802 578952
rect 213177 578370 213243 578373
rect 210742 578368 213243 578370
rect 210742 578312 213182 578368
rect 213238 578312 213243 578368
rect 210742 578310 213243 578312
rect 300718 578370 300778 578952
rect 302325 578370 302391 578373
rect 300718 578368 302391 578370
rect 300718 578312 302330 578368
rect 302386 578312 302391 578368
rect 300718 578310 302391 578312
rect 213177 578307 213243 578310
rect 302325 578307 302391 578310
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 583520 577540 584960 577630
rect 58525 576874 58591 576877
rect 59494 576874 60076 576910
rect 58525 576872 60076 576874
rect 58525 576816 58530 576872
rect 58586 576850 60076 576872
rect 147029 576874 147095 576877
rect 149470 576874 150052 576910
rect 147029 576872 150052 576874
rect 58586 576816 59554 576850
rect 58525 576814 59554 576816
rect 147029 576816 147034 576872
rect 147090 576850 150052 576872
rect 237373 576874 237439 576877
rect 239446 576874 240120 576910
rect 237373 576872 240120 576874
rect 147090 576816 149530 576850
rect 147029 576814 149530 576816
rect 237373 576816 237378 576872
rect 237434 576850 240120 576872
rect 237434 576816 239506 576850
rect 237373 576814 239506 576816
rect 58525 576811 58591 576814
rect 147029 576811 147095 576814
rect 237373 576811 237439 576814
rect 120766 575650 120826 576232
rect 210742 575653 210802 576232
rect 123477 575650 123543 575653
rect 120766 575648 123543 575650
rect 120766 575592 123482 575648
rect 123538 575592 123543 575648
rect 120766 575590 123543 575592
rect 210742 575648 210851 575653
rect 210742 575592 210790 575648
rect 210846 575592 210851 575648
rect 210742 575590 210851 575592
rect 300718 575650 300778 576232
rect 301589 575650 301655 575653
rect 300718 575648 301655 575650
rect 300718 575592 301594 575648
rect 301650 575592 301655 575648
rect 300718 575590 301655 575592
rect 123477 575587 123543 575590
rect 210785 575587 210851 575590
rect 301589 575587 301655 575590
rect 433382 574565 433442 575076
rect 433382 574560 433491 574565
rect 433382 574504 433430 574560
rect 433486 574504 433491 574560
rect 433382 574502 433491 574504
rect 433425 574499 433491 574502
rect 321553 574426 321619 574429
rect 321553 574424 325036 574426
rect 321553 574368 321558 574424
rect 321614 574368 325036 574424
rect 321553 574366 325036 574368
rect 321553 574363 321619 574366
rect 57789 573474 57855 573477
rect 59494 573474 60076 573510
rect 57789 573472 60076 573474
rect 57789 573416 57794 573472
rect 57850 573450 60076 573472
rect 149053 573474 149119 573477
rect 149470 573474 150052 573510
rect 149053 573472 150052 573474
rect 57850 573416 59554 573450
rect 57789 573414 59554 573416
rect 149053 573416 149058 573472
rect 149114 573450 150052 573472
rect 237373 573474 237439 573477
rect 239446 573474 240120 573510
rect 237373 573472 240120 573474
rect 149114 573416 149530 573450
rect 149053 573414 149530 573416
rect 237373 573416 237378 573472
rect 237434 573450 240120 573472
rect 237434 573416 239506 573450
rect 237373 573414 239506 573416
rect 57789 573411 57855 573414
rect 149053 573411 149119 573414
rect 237373 573411 237439 573414
rect 120766 572794 120826 572832
rect 122281 572794 122347 572797
rect 120766 572792 122347 572794
rect 120766 572736 122286 572792
rect 122342 572736 122347 572792
rect 120766 572734 122347 572736
rect 210742 572794 210802 572832
rect 213361 572794 213427 572797
rect 210742 572792 213427 572794
rect 210742 572736 213366 572792
rect 213422 572736 213427 572792
rect 210742 572734 213427 572736
rect 300718 572794 300778 572832
rect 303061 572794 303127 572797
rect 300718 572792 303127 572794
rect 300718 572736 303066 572792
rect 303122 572736 303127 572792
rect 300718 572734 303127 572736
rect 122281 572731 122347 572734
rect 213361 572731 213427 572734
rect 303061 572731 303127 572734
rect 59537 570790 59603 570793
rect 59537 570788 60076 570790
rect 59537 570732 59542 570788
rect 59598 570732 60076 570788
rect 59537 570730 60076 570732
rect 148225 570754 148291 570757
rect 149470 570754 150052 570790
rect 148225 570752 150052 570754
rect 59537 570727 59603 570730
rect 148225 570696 148230 570752
rect 148286 570730 150052 570752
rect 237373 570754 237439 570757
rect 239446 570754 240120 570790
rect 237373 570752 240120 570754
rect 148286 570696 149530 570730
rect 148225 570694 149530 570696
rect 237373 570696 237378 570752
rect 237434 570730 240120 570752
rect 237434 570696 239506 570730
rect 237373 570694 239506 570696
rect 148225 570691 148291 570694
rect 237373 570691 237439 570694
rect 210877 570346 210943 570349
rect 436369 570346 436435 570349
rect 210742 570344 210943 570346
rect 210742 570288 210882 570344
rect 210938 570288 210943 570344
rect 210742 570286 210943 570288
rect 433780 570344 436435 570346
rect 433780 570288 436374 570344
rect 436430 570288 436435 570344
rect 433780 570286 436435 570288
rect 210742 570112 210802 570286
rect 210877 570283 210943 570286
rect 436369 570283 436435 570286
rect 120766 570074 120826 570112
rect 121545 570074 121611 570077
rect 120766 570072 121611 570074
rect 120766 570016 121550 570072
rect 121606 570016 121611 570072
rect 120766 570014 121611 570016
rect 300718 570074 300778 570112
rect 301681 570074 301747 570077
rect 300718 570072 301747 570074
rect 300718 570016 301686 570072
rect 301742 570016 301747 570072
rect 300718 570014 301747 570016
rect 121545 570011 121611 570014
rect 301681 570011 301747 570014
rect 321553 569666 321619 569669
rect 321553 569664 325036 569666
rect 321553 569608 321558 569664
rect 321614 569608 325036 569664
rect 321553 569606 325036 569608
rect 321553 569603 321619 569606
rect -960 566796 480 567036
rect 436461 565586 436527 565589
rect 433780 565584 436527 565586
rect 433780 565528 436466 565584
rect 436522 565528 436527 565584
rect 433780 565526 436527 565528
rect 436461 565523 436527 565526
rect 321553 564906 321619 564909
rect 321553 564904 325036 564906
rect 321553 564848 321558 564904
rect 321614 564848 325036 564904
rect 321553 564846 325036 564848
rect 321553 564843 321619 564846
rect 583520 564212 584960 564452
rect 433566 560421 433626 560796
rect 433517 560416 433626 560421
rect 433517 560360 433522 560416
rect 433578 560360 433626 560416
rect 433517 560358 433626 560360
rect 433517 560355 433583 560358
rect 321553 560146 321619 560149
rect 321553 560144 325036 560146
rect 321553 560088 321558 560144
rect 321614 560088 325036 560144
rect 321553 560086 325036 560088
rect 321553 560083 321619 560086
rect 436553 556066 436619 556069
rect 433780 556064 436619 556066
rect 433780 556008 436558 556064
rect 436614 556008 436619 556064
rect 433780 556006 436619 556008
rect 436553 556003 436619 556006
rect 321553 555386 321619 555389
rect 321553 555384 325036 555386
rect 321553 555328 321558 555384
rect 321614 555328 325036 555384
rect 321553 555326 325036 555328
rect 321553 555323 321619 555326
rect -960 553740 480 553980
rect 68093 552666 68159 552669
rect 121678 552666 121684 552668
rect 68093 552664 121684 552666
rect 68093 552608 68098 552664
rect 68154 552608 121684 552664
rect 68093 552606 121684 552608
rect 68093 552603 68159 552606
rect 121678 552604 121684 552606
rect 121748 552604 121754 552668
rect 436645 551306 436711 551309
rect 433780 551304 436711 551306
rect 433780 551248 436650 551304
rect 436706 551248 436711 551304
rect 433780 551246 436711 551248
rect 436645 551243 436711 551246
rect 583520 551020 584960 551260
rect 320817 550626 320883 550629
rect 320817 550624 325036 550626
rect 320817 550568 320822 550624
rect 320878 550568 325036 550624
rect 320817 550566 325036 550568
rect 320817 550563 320883 550566
rect 298093 550218 298159 550221
rect 320909 550218 320975 550221
rect 298093 550216 320975 550218
rect 298093 550160 298098 550216
rect 298154 550160 320914 550216
rect 320970 550160 320975 550216
rect 298093 550158 320975 550160
rect 298093 550155 298159 550158
rect 320909 550155 320975 550158
rect 297357 550082 297423 550085
rect 322197 550082 322263 550085
rect 297357 550080 322263 550082
rect 297357 550024 297362 550080
rect 297418 550024 322202 550080
rect 322258 550024 322263 550080
rect 297357 550022 322263 550024
rect 297357 550019 297423 550022
rect 322197 550019 322263 550022
rect 245837 549946 245903 549949
rect 323669 549946 323735 549949
rect 245837 549944 323735 549946
rect 245837 549888 245842 549944
rect 245898 549888 323674 549944
rect 323730 549888 323735 549944
rect 245837 549886 323735 549888
rect 245837 549883 245903 549886
rect 323669 549883 323735 549886
rect 248689 549810 248755 549813
rect 301773 549810 301839 549813
rect 248689 549808 301839 549810
rect 248689 549752 248694 549808
rect 248750 549752 301778 549808
rect 301834 549752 301839 549808
rect 248689 549750 301839 549752
rect 248689 549747 248755 549750
rect 301773 549747 301839 549750
rect 241513 549674 241579 549677
rect 301957 549674 302023 549677
rect 241513 549672 302023 549674
rect 241513 549616 241518 549672
rect 241574 549616 301962 549672
rect 302018 549616 302023 549672
rect 241513 549614 302023 549616
rect 241513 549611 241579 549614
rect 301957 549611 302023 549614
rect 238661 549538 238727 549541
rect 299974 549538 299980 549540
rect 238661 549536 299980 549538
rect 238661 549480 238666 549536
rect 238722 549480 299980 549536
rect 238661 549478 299980 549480
rect 238661 549475 238727 549478
rect 299974 549476 299980 549478
rect 300044 549476 300050 549540
rect 255129 549402 255195 549405
rect 321093 549402 321159 549405
rect 255129 549400 321159 549402
rect 255129 549344 255134 549400
rect 255190 549344 321098 549400
rect 321154 549344 321159 549400
rect 255129 549342 321159 549344
rect 255129 549339 255195 549342
rect 321093 549339 321159 549342
rect 237189 548178 237255 548181
rect 293769 548178 293835 548181
rect 237189 548176 238770 548178
rect 237189 548120 237194 548176
rect 237250 548120 238770 548176
rect 237189 548118 238770 548120
rect 237189 548115 237255 548118
rect 238710 547906 238770 548118
rect 293769 548176 296730 548178
rect 293769 548120 293774 548176
rect 293830 548120 296730 548176
rect 293769 548118 296730 548120
rect 293769 548115 293835 548118
rect 296670 548042 296730 548118
rect 317229 548042 317295 548045
rect 296670 548040 317295 548042
rect 296670 547984 317234 548040
rect 317290 547984 317295 548040
rect 296670 547982 317295 547984
rect 317229 547979 317295 547982
rect 301865 547906 301931 547909
rect 238710 547904 301931 547906
rect 238710 547848 301870 547904
rect 301926 547848 301931 547904
rect 238710 547846 301931 547848
rect 301865 547843 301931 547846
rect 433566 546413 433626 546516
rect 433566 546408 433675 546413
rect 433566 546352 433614 546408
rect 433670 546352 433675 546408
rect 433566 546350 433675 546352
rect 433609 546347 433675 546350
rect 321829 545866 321895 545869
rect 321829 545864 325036 545866
rect 321829 545808 321834 545864
rect 321890 545808 325036 545864
rect 321829 545806 325036 545808
rect 321829 545803 321895 545806
rect 436737 541786 436803 541789
rect 433780 541784 436803 541786
rect 433780 541728 436742 541784
rect 436798 541728 436803 541784
rect 433780 541726 436803 541728
rect 436737 541723 436803 541726
rect 321553 541106 321619 541109
rect 321553 541104 325036 541106
rect 321553 541048 321558 541104
rect 321614 541048 325036 541104
rect 321553 541046 325036 541048
rect 321553 541043 321619 541046
rect -960 540684 480 540924
rect 302601 540426 302667 540429
rect 299828 540424 302667 540426
rect 299828 540368 302606 540424
rect 302662 540368 302667 540424
rect 299828 540366 302667 540368
rect 302601 540363 302667 540366
rect 583520 537692 584960 537932
rect 436185 537026 436251 537029
rect 433780 537024 436251 537026
rect 433780 536968 436190 537024
rect 436246 536968 436251 537024
rect 433780 536966 436251 536968
rect 436185 536963 436251 536966
rect 321553 536346 321619 536349
rect 321553 536344 325036 536346
rect 321553 536288 321558 536344
rect 321614 536288 325036 536344
rect 321553 536286 325036 536288
rect 321553 536283 321619 536286
rect 434805 532266 434871 532269
rect 433780 532264 434871 532266
rect 433780 532208 434810 532264
rect 434866 532208 434871 532264
rect 433780 532206 434871 532208
rect 434805 532203 434871 532206
rect 322197 531586 322263 531589
rect 322197 531584 325036 531586
rect 322197 531528 322202 531584
rect 322258 531528 325036 531584
rect 322197 531526 325036 531528
rect 322197 531523 322263 531526
rect -960 527764 480 528004
rect 436277 527506 436343 527509
rect 433780 527504 436343 527506
rect 433780 527448 436282 527504
rect 436338 527448 436343 527504
rect 433780 527446 436343 527448
rect 436277 527443 436343 527446
rect 321553 526826 321619 526829
rect 321553 526824 325036 526826
rect 321553 526768 321558 526824
rect 321614 526768 325036 526824
rect 321553 526766 325036 526768
rect 321553 526763 321619 526766
rect 302969 525466 303035 525469
rect 299828 525464 303035 525466
rect 299828 525408 302974 525464
rect 303030 525408 303035 525464
rect 299828 525406 303035 525408
rect 302969 525403 303035 525406
rect 583520 524364 584960 524604
rect 433566 522613 433626 522716
rect 299974 522548 299980 522612
rect 300044 522610 300050 522612
rect 300044 522550 433258 522610
rect 300044 522548 300050 522550
rect 301957 522474 302023 522477
rect 433198 522474 433258 522550
rect 433517 522608 433626 522613
rect 433517 522552 433522 522608
rect 433578 522552 433626 522608
rect 433517 522550 433626 522552
rect 433517 522547 433583 522550
rect 436369 522474 436435 522477
rect 301957 522472 431970 522474
rect 301957 522416 301962 522472
rect 302018 522416 431970 522472
rect 301957 522414 431970 522416
rect 433198 522472 436435 522474
rect 433198 522416 436374 522472
rect 436430 522416 436435 522472
rect 433198 522414 436435 522416
rect 301957 522411 302023 522414
rect 431910 522338 431970 522414
rect 436369 522411 436435 522414
rect 436134 522338 436140 522340
rect 431910 522278 436140 522338
rect 436134 522276 436140 522278
rect 436204 522276 436210 522340
rect 301497 520162 301563 520165
rect 429193 520162 429259 520165
rect 301497 520160 429259 520162
rect 301497 520104 301502 520160
rect 301558 520104 429198 520160
rect 429254 520104 429259 520160
rect 301497 520102 429259 520104
rect 301497 520099 301563 520102
rect 429193 520099 429259 520102
rect 329741 520026 329807 520029
rect 434713 520026 434779 520029
rect 329741 520024 434779 520026
rect 329741 519968 329746 520024
rect 329802 519968 434718 520024
rect 434774 519968 434779 520024
rect 329741 519966 434779 519968
rect 329741 519963 329807 519966
rect 434713 519963 434779 519966
rect 57881 517986 57947 517989
rect 57881 517984 60076 517986
rect 57881 517928 57886 517984
rect 57942 517928 60076 517984
rect 57881 517926 60076 517928
rect 57881 517923 57947 517926
rect 360878 516700 360884 516764
rect 360948 516762 360954 516764
rect 397453 516762 397519 516765
rect 360948 516760 397519 516762
rect 360948 516704 397458 516760
rect 397514 516704 397519 516760
rect 360948 516702 397519 516704
rect 360948 516700 360954 516702
rect 397453 516699 397519 516702
rect 363454 515340 363460 515404
rect 363524 515402 363530 515404
rect 506473 515402 506539 515405
rect 363524 515400 506539 515402
rect 363524 515344 506478 515400
rect 506534 515344 506539 515400
rect 363524 515342 506539 515344
rect 363524 515340 363530 515342
rect 506473 515339 506539 515342
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 302693 510506 302759 510509
rect 299828 510504 302759 510506
rect 299828 510448 302698 510504
rect 302754 510448 302759 510504
rect 299828 510446 302759 510448
rect 302693 510443 302759 510446
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect 302233 495546 302299 495549
rect 299828 495544 302299 495546
rect 299828 495488 302238 495544
rect 302294 495488 302299 495544
rect 299828 495486 302299 495488
rect 302233 495483 302299 495486
rect 363638 491812 363644 491876
rect 363708 491874 363714 491876
rect 476062 491874 476068 491876
rect 363708 491814 476068 491874
rect 363708 491812 363714 491814
rect 476062 491812 476068 491814
rect 476132 491812 476138 491876
rect 367686 490452 367692 490516
rect 367756 490514 367762 490516
rect 483013 490514 483079 490517
rect 367756 490512 483079 490514
rect 367756 490456 483018 490512
rect 483074 490456 483079 490512
rect 367756 490454 483079 490456
rect 367756 490452 367762 490454
rect 483013 490451 483079 490454
rect -960 488596 480 488836
rect 367870 487732 367876 487796
rect 367940 487794 367946 487796
rect 511993 487794 512059 487797
rect 367940 487792 512059 487794
rect 367940 487736 511998 487792
rect 512054 487736 512059 487792
rect 367940 487734 512059 487736
rect 367940 487732 367946 487734
rect 511993 487731 512059 487734
rect 206134 486372 206140 486436
rect 206204 486434 206210 486436
rect 488574 486434 488580 486436
rect 206204 486374 488580 486434
rect 206204 486372 206210 486374
rect 488574 486372 488580 486374
rect 488644 486372 488650 486436
rect 59302 485692 59308 485756
rect 59372 485754 59378 485756
rect 72509 485754 72575 485757
rect 59372 485752 72575 485754
rect 59372 485696 72514 485752
rect 72570 485696 72575 485752
rect 59372 485694 72575 485696
rect 59372 485692 59378 485694
rect 72509 485691 72575 485694
rect 158621 485754 158687 485757
rect 182265 485754 182331 485757
rect 158621 485752 182331 485754
rect 158621 485696 158626 485752
rect 158682 485696 182270 485752
rect 182326 485696 182331 485752
rect 158621 485694 182331 485696
rect 158621 485691 158687 485694
rect 182265 485691 182331 485694
rect 184841 485754 184907 485757
rect 196750 485754 196756 485756
rect 184841 485752 196756 485754
rect 184841 485696 184846 485752
rect 184902 485696 196756 485752
rect 184841 485694 196756 485696
rect 184841 485691 184907 485694
rect 196750 485692 196756 485694
rect 196820 485692 196826 485756
rect 211153 485754 211219 485757
rect 212390 485754 212396 485756
rect 211153 485752 212396 485754
rect 211153 485696 211158 485752
rect 211214 485696 212396 485752
rect 211153 485694 212396 485696
rect 211153 485691 211219 485694
rect 212390 485692 212396 485694
rect 212460 485692 212466 485756
rect 235809 485754 235875 485757
rect 357934 485754 357940 485756
rect 235809 485752 357940 485754
rect 235809 485696 235814 485752
rect 235870 485696 357940 485752
rect 235809 485694 357940 485696
rect 235809 485691 235875 485694
rect 357934 485692 357940 485694
rect 358004 485692 358010 485756
rect 54702 485556 54708 485620
rect 54772 485618 54778 485620
rect 73797 485618 73863 485621
rect 54772 485616 73863 485618
rect 54772 485560 73802 485616
rect 73858 485560 73863 485616
rect 54772 485558 73863 485560
rect 54772 485556 54778 485558
rect 73797 485555 73863 485558
rect 171133 485618 171199 485621
rect 202270 485618 202276 485620
rect 171133 485616 202276 485618
rect 171133 485560 171138 485616
rect 171194 485560 202276 485616
rect 171133 485558 202276 485560
rect 171133 485555 171199 485558
rect 202270 485556 202276 485558
rect 202340 485556 202346 485620
rect 212533 485618 212599 485621
rect 213678 485618 213684 485620
rect 212533 485616 213684 485618
rect 212533 485560 212538 485616
rect 212594 485560 213684 485616
rect 212533 485558 213684 485560
rect 212533 485555 212599 485558
rect 213678 485556 213684 485558
rect 213748 485556 213754 485620
rect 230657 485618 230723 485621
rect 364926 485618 364932 485620
rect 230657 485616 364932 485618
rect 230657 485560 230662 485616
rect 230718 485560 364932 485616
rect 230657 485558 364932 485560
rect 230657 485555 230723 485558
rect 364926 485556 364932 485558
rect 364996 485556 365002 485620
rect 51942 485420 51948 485484
rect 52012 485482 52018 485484
rect 74257 485482 74323 485485
rect 52012 485480 74323 485482
rect 52012 485424 74262 485480
rect 74318 485424 74323 485480
rect 52012 485422 74323 485424
rect 52012 485420 52018 485422
rect 74257 485419 74323 485422
rect 74441 485482 74507 485485
rect 79961 485482 80027 485485
rect 74441 485480 80027 485482
rect 74441 485424 74446 485480
rect 74502 485424 79966 485480
rect 80022 485424 80027 485480
rect 74441 485422 80027 485424
rect 74441 485419 74507 485422
rect 79961 485419 80027 485422
rect 163681 485482 163747 485485
rect 196566 485482 196572 485484
rect 163681 485480 196572 485482
rect 163681 485424 163686 485480
rect 163742 485424 196572 485480
rect 163681 485422 196572 485424
rect 163681 485419 163747 485422
rect 196566 485420 196572 485422
rect 196636 485420 196642 485484
rect 234337 485482 234403 485485
rect 371734 485482 371740 485484
rect 234337 485480 371740 485482
rect 234337 485424 234342 485480
rect 234398 485424 371740 485480
rect 234337 485422 371740 485424
rect 234337 485419 234403 485422
rect 371734 485420 371740 485422
rect 371804 485420 371810 485484
rect 53414 485284 53420 485348
rect 53484 485346 53490 485348
rect 76005 485346 76071 485349
rect 53484 485344 76071 485346
rect 53484 485288 76010 485344
rect 76066 485288 76071 485344
rect 53484 485286 76071 485288
rect 53484 485284 53490 485286
rect 76005 485283 76071 485286
rect 145649 485346 145715 485349
rect 197854 485346 197860 485348
rect 145649 485344 197860 485346
rect 145649 485288 145654 485344
rect 145710 485288 197860 485344
rect 145649 485286 197860 485288
rect 145649 485283 145715 485286
rect 197854 485284 197860 485286
rect 197924 485284 197930 485348
rect 200205 485346 200271 485349
rect 217542 485346 217548 485348
rect 200205 485344 217548 485346
rect 200205 485288 200210 485344
rect 200266 485288 217548 485344
rect 200205 485286 217548 485288
rect 200205 485283 200271 485286
rect 217542 485284 217548 485286
rect 217612 485284 217618 485348
rect 235901 485346 235967 485349
rect 373758 485346 373764 485348
rect 235901 485344 373764 485346
rect 235901 485288 235906 485344
rect 235962 485288 373764 485344
rect 235901 485286 373764 485288
rect 235901 485283 235967 485286
rect 373758 485284 373764 485286
rect 373828 485284 373834 485348
rect 50286 485148 50292 485212
rect 50356 485210 50362 485212
rect 77293 485210 77359 485213
rect 50356 485208 77359 485210
rect 50356 485152 77298 485208
rect 77354 485152 77359 485208
rect 50356 485150 77359 485152
rect 50356 485148 50362 485150
rect 77293 485147 77359 485150
rect 147581 485210 147647 485213
rect 191097 485210 191163 485213
rect 147581 485208 191163 485210
rect 147581 485152 147586 485208
rect 147642 485152 191102 485208
rect 191158 485152 191163 485208
rect 147581 485150 191163 485152
rect 147581 485147 147647 485150
rect 191097 485147 191163 485150
rect 197353 485210 197419 485213
rect 198590 485210 198596 485212
rect 197353 485208 198596 485210
rect 197353 485152 197358 485208
rect 197414 485152 198596 485208
rect 197353 485150 198596 485152
rect 197353 485147 197419 485150
rect 198590 485148 198596 485150
rect 198660 485148 198666 485212
rect 204437 485210 204503 485213
rect 205398 485210 205404 485212
rect 204437 485208 205404 485210
rect 204437 485152 204442 485208
rect 204498 485152 205404 485208
rect 204437 485150 205404 485152
rect 204437 485147 204503 485150
rect 205398 485148 205404 485150
rect 205468 485148 205474 485212
rect 206185 485210 206251 485213
rect 206870 485210 206876 485212
rect 206185 485208 206876 485210
rect 206185 485152 206190 485208
rect 206246 485152 206876 485208
rect 206185 485150 206876 485152
rect 206185 485147 206251 485150
rect 206870 485148 206876 485150
rect 206940 485148 206946 485212
rect 219198 485148 219204 485212
rect 219268 485210 219274 485212
rect 225689 485210 225755 485213
rect 219268 485208 225755 485210
rect 219268 485152 225694 485208
rect 225750 485152 225755 485208
rect 219268 485150 225755 485152
rect 219268 485148 219274 485150
rect 225689 485147 225755 485150
rect 232313 485210 232379 485213
rect 374494 485210 374500 485212
rect 232313 485208 374500 485210
rect 232313 485152 232318 485208
rect 232374 485152 374500 485208
rect 232313 485150 374500 485152
rect 232313 485147 232379 485150
rect 374494 485148 374500 485150
rect 374564 485148 374570 485212
rect 57830 485012 57836 485076
rect 57900 485074 57906 485076
rect 91369 485074 91435 485077
rect 57900 485072 91435 485074
rect 57900 485016 91374 485072
rect 91430 485016 91435 485072
rect 57900 485014 91435 485016
rect 57900 485012 57906 485014
rect 91369 485011 91435 485014
rect 145465 485074 145531 485077
rect 200614 485074 200620 485076
rect 145465 485072 200620 485074
rect 145465 485016 145470 485072
rect 145526 485016 200620 485072
rect 145465 485014 200620 485016
rect 145465 485011 145531 485014
rect 200614 485012 200620 485014
rect 200684 485012 200690 485076
rect 208393 485074 208459 485077
rect 208894 485074 208900 485076
rect 208393 485072 208900 485074
rect 208393 485016 208398 485072
rect 208454 485016 208900 485072
rect 208393 485014 208900 485016
rect 208393 485011 208459 485014
rect 208894 485012 208900 485014
rect 208964 485012 208970 485076
rect 219014 485012 219020 485076
rect 219084 485074 219090 485076
rect 226149 485074 226215 485077
rect 219084 485072 226215 485074
rect 219084 485016 226154 485072
rect 226210 485016 226215 485072
rect 219084 485014 226215 485016
rect 219084 485012 219090 485014
rect 226149 485011 226215 485014
rect 231761 485074 231827 485077
rect 375966 485074 375972 485076
rect 231761 485072 375972 485074
rect 231761 485016 231766 485072
rect 231822 485016 375972 485072
rect 231761 485014 375972 485016
rect 231761 485011 231827 485014
rect 375966 485012 375972 485014
rect 376036 485012 376042 485076
rect 59118 484876 59124 484940
rect 59188 484938 59194 484940
rect 68921 484938 68987 484941
rect 59188 484936 68987 484938
rect 59188 484880 68926 484936
rect 68982 484880 68987 484936
rect 59188 484878 68987 484880
rect 59188 484876 59194 484878
rect 68921 484875 68987 484878
rect 187049 484938 187115 484941
rect 198038 484938 198044 484940
rect 187049 484936 198044 484938
rect 187049 484880 187054 484936
rect 187110 484880 198044 484936
rect 187049 484878 198044 484880
rect 187049 484875 187115 484878
rect 198038 484876 198044 484878
rect 198108 484876 198114 484940
rect 201493 484938 201559 484941
rect 202638 484938 202644 484940
rect 201493 484936 202644 484938
rect 201493 484880 201498 484936
rect 201554 484880 202644 484936
rect 201493 484878 202644 484880
rect 201493 484875 201559 484878
rect 202638 484876 202644 484878
rect 202708 484876 202714 484940
rect 248689 484938 248755 484941
rect 356646 484938 356652 484940
rect 248689 484936 356652 484938
rect 248689 484880 248694 484936
rect 248750 484880 356652 484936
rect 248689 484878 356652 484880
rect 248689 484875 248755 484878
rect 356646 484876 356652 484878
rect 356716 484876 356722 484940
rect 197353 484802 197419 484805
rect 198406 484802 198412 484804
rect 197353 484800 198412 484802
rect 197353 484744 197358 484800
rect 197414 484744 198412 484800
rect 197353 484742 198412 484744
rect 197353 484739 197419 484742
rect 198406 484740 198412 484742
rect 198476 484740 198482 484804
rect 200481 484802 200547 484805
rect 201350 484802 201356 484804
rect 200481 484800 201356 484802
rect 200481 484744 200486 484800
rect 200542 484744 201356 484800
rect 200481 484742 201356 484744
rect 200481 484739 200547 484742
rect 201350 484740 201356 484742
rect 201420 484740 201426 484804
rect 208393 484802 208459 484805
rect 209078 484802 209084 484804
rect 208393 484800 209084 484802
rect 208393 484744 208398 484800
rect 208454 484744 209084 484800
rect 208393 484742 209084 484744
rect 208393 484739 208459 484742
rect 209078 484740 209084 484742
rect 209148 484740 209154 484804
rect 191097 484666 191163 484669
rect 200798 484666 200804 484668
rect 191097 484664 200804 484666
rect 191097 484608 191102 484664
rect 191158 484608 200804 484664
rect 191097 484606 200804 484608
rect 191097 484603 191163 484606
rect 200798 484604 200804 484606
rect 200868 484604 200874 484668
rect 211153 484666 211219 484669
rect 211654 484666 211660 484668
rect 211153 484664 211660 484666
rect 211153 484608 211158 484664
rect 211214 484608 211660 484664
rect 211153 484606 211660 484608
rect 211153 484603 211219 484606
rect 211654 484604 211660 484606
rect 211724 484604 211730 484668
rect 53281 484532 53347 484533
rect 53649 484532 53715 484533
rect 53230 484530 53236 484532
rect 53190 484470 53236 484530
rect 53300 484528 53347 484532
rect 53598 484530 53604 484532
rect 53342 484472 53347 484528
rect 53230 484468 53236 484470
rect 53300 484468 53347 484472
rect 53558 484470 53604 484530
rect 53668 484528 53715 484532
rect 53710 484472 53715 484528
rect 53598 484468 53604 484470
rect 53668 484468 53715 484472
rect 53281 484467 53347 484468
rect 53649 484467 53715 484468
rect 214741 484530 214807 484533
rect 216990 484530 216996 484532
rect 214741 484528 216996 484530
rect 214741 484472 214746 484528
rect 214802 484472 216996 484528
rect 214741 484470 216996 484472
rect 214741 484467 214807 484470
rect 216990 484468 216996 484470
rect 217060 484468 217066 484532
rect 219934 484468 219940 484532
rect 220004 484530 220010 484532
rect 224861 484530 224927 484533
rect 220004 484528 224927 484530
rect 220004 484472 224866 484528
rect 224922 484472 224927 484528
rect 583520 484516 584960 484756
rect 220004 484470 224927 484472
rect 220004 484468 220010 484470
rect 224861 484467 224927 484470
rect 281073 483986 281139 483989
rect 377438 483986 377444 483988
rect 281073 483984 377444 483986
rect 281073 483928 281078 483984
rect 281134 483928 377444 483984
rect 281073 483926 377444 483928
rect 281073 483923 281139 483926
rect 377438 483924 377444 483926
rect 377508 483924 377514 483988
rect 156505 483850 156571 483853
rect 205766 483850 205772 483852
rect 156505 483848 205772 483850
rect 156505 483792 156510 483848
rect 156566 483792 205772 483848
rect 156505 483790 205772 483792
rect 156505 483787 156571 483790
rect 205766 483788 205772 483790
rect 205836 483788 205842 483852
rect 252921 483850 252987 483853
rect 377254 483850 377260 483852
rect 252921 483848 377260 483850
rect 252921 483792 252926 483848
rect 252982 483792 377260 483848
rect 252921 483790 377260 483792
rect 252921 483787 252987 483790
rect 377254 483788 377260 483790
rect 377324 483788 377330 483852
rect 150249 483714 150315 483717
rect 213126 483714 213132 483716
rect 150249 483712 213132 483714
rect 150249 483656 150254 483712
rect 150310 483656 213132 483712
rect 150249 483654 213132 483656
rect 150249 483651 150315 483654
rect 213126 483652 213132 483654
rect 213196 483652 213202 483716
rect 230381 483714 230447 483717
rect 360694 483714 360700 483716
rect 230381 483712 360700 483714
rect 230381 483656 230386 483712
rect 230442 483656 360700 483712
rect 230381 483654 360700 483656
rect 230381 483651 230447 483654
rect 360694 483652 360700 483654
rect 360764 483652 360770 483716
rect 46790 482836 46796 482900
rect 46860 482898 46866 482900
rect 66345 482898 66411 482901
rect 46860 482896 66411 482898
rect 46860 482840 66350 482896
rect 66406 482840 66411 482896
rect 46860 482838 66411 482840
rect 46860 482836 46866 482838
rect 66345 482835 66411 482838
rect 47710 482700 47716 482764
rect 47780 482762 47786 482764
rect 120441 482762 120507 482765
rect 47780 482760 120507 482762
rect 47780 482704 120446 482760
rect 120502 482704 120507 482760
rect 47780 482702 120507 482704
rect 47780 482700 47786 482702
rect 120441 482699 120507 482702
rect 46565 482626 46631 482629
rect 120901 482626 120967 482629
rect 46565 482624 120967 482626
rect 46565 482568 46570 482624
rect 46626 482568 120906 482624
rect 120962 482568 120967 482624
rect 46565 482566 120967 482568
rect 46565 482563 46631 482566
rect 120901 482563 120967 482566
rect 46473 482490 46539 482493
rect 120073 482490 120139 482493
rect 46473 482488 120139 482490
rect 46473 482432 46478 482488
rect 46534 482432 120078 482488
rect 120134 482432 120139 482488
rect 46473 482430 120139 482432
rect 46473 482427 46539 482430
rect 120073 482427 120139 482430
rect 236361 482490 236427 482493
rect 375414 482490 375420 482492
rect 236361 482488 375420 482490
rect 236361 482432 236366 482488
rect 236422 482432 375420 482488
rect 236361 482430 375420 482432
rect 236361 482427 236427 482430
rect 375414 482428 375420 482430
rect 375484 482428 375490 482492
rect 43897 482354 43963 482357
rect 121361 482354 121427 482357
rect 43897 482352 121427 482354
rect 43897 482296 43902 482352
rect 43958 482296 121366 482352
rect 121422 482296 121427 482352
rect 43897 482294 121427 482296
rect 43897 482291 43963 482294
rect 121361 482291 121427 482294
rect 155861 482354 155927 482357
rect 213862 482354 213868 482356
rect 155861 482352 213868 482354
rect 155861 482296 155866 482352
rect 155922 482296 213868 482352
rect 155861 482294 213868 482296
rect 155861 482291 155927 482294
rect 213862 482292 213868 482294
rect 213932 482292 213938 482356
rect 222561 482354 222627 482357
rect 376150 482354 376156 482356
rect 222561 482352 376156 482354
rect 222561 482296 222566 482352
rect 222622 482296 376156 482352
rect 222561 482294 376156 482296
rect 222561 482291 222627 482294
rect 376150 482292 376156 482294
rect 376220 482292 376226 482356
rect 3417 482218 3483 482221
rect 316677 482218 316743 482221
rect 3417 482216 316743 482218
rect 3417 482160 3422 482216
rect 3478 482160 316682 482216
rect 316738 482160 316743 482216
rect 3417 482158 316743 482160
rect 3417 482155 3483 482158
rect 316677 482155 316743 482158
rect 155217 480994 155283 480997
rect 215334 480994 215340 480996
rect 155217 480992 215340 480994
rect 155217 480936 155222 480992
rect 155278 480936 215340 480992
rect 155217 480934 215340 480936
rect 155217 480931 155283 480934
rect 215334 480932 215340 480934
rect 215404 480932 215410 480996
rect 247309 480994 247375 480997
rect 374862 480994 374868 480996
rect 247309 480992 374868 480994
rect 247309 480936 247314 480992
rect 247370 480936 374868 480992
rect 247309 480934 374868 480936
rect 247309 480931 247375 480934
rect 374862 480932 374868 480934
rect 374932 480932 374938 480996
rect 147213 480858 147279 480861
rect 215886 480858 215892 480860
rect 147213 480856 215892 480858
rect 147213 480800 147218 480856
rect 147274 480800 215892 480856
rect 147213 480798 215892 480800
rect 147213 480795 147279 480798
rect 215886 480796 215892 480798
rect 215956 480796 215962 480860
rect 232129 480858 232195 480861
rect 370078 480858 370084 480860
rect 232129 480856 370084 480858
rect 232129 480800 232134 480856
rect 232190 480800 370084 480856
rect 232129 480798 370084 480800
rect 232129 480795 232195 480798
rect 370078 480796 370084 480798
rect 370148 480796 370154 480860
rect 42609 480042 42675 480045
rect 80513 480042 80579 480045
rect 42609 480040 80579 480042
rect 42609 479984 42614 480040
rect 42670 479984 80518 480040
rect 80574 479984 80579 480040
rect 42609 479982 80579 479984
rect 42609 479979 42675 479982
rect 80513 479979 80579 479982
rect 57462 479844 57468 479908
rect 57532 479906 57538 479908
rect 118785 479906 118851 479909
rect 57532 479904 118851 479906
rect 57532 479848 118790 479904
rect 118846 479848 118851 479904
rect 57532 479846 118851 479848
rect 57532 479844 57538 479846
rect 118785 479843 118851 479846
rect 57094 479708 57100 479772
rect 57164 479770 57170 479772
rect 122373 479770 122439 479773
rect 57164 479768 122439 479770
rect 57164 479712 122378 479768
rect 122434 479712 122439 479768
rect 57164 479710 122439 479712
rect 57164 479708 57170 479710
rect 122373 479707 122439 479710
rect 178677 479770 178743 479773
rect 217174 479770 217180 479772
rect 178677 479768 217180 479770
rect 178677 479712 178682 479768
rect 178738 479712 217180 479768
rect 178677 479710 217180 479712
rect 178677 479707 178743 479710
rect 217174 479708 217180 479710
rect 217244 479708 217250 479772
rect 44950 479572 44956 479636
rect 45020 479634 45026 479636
rect 117957 479634 118023 479637
rect 45020 479632 118023 479634
rect 45020 479576 117962 479632
rect 118018 479576 118023 479632
rect 45020 479574 118023 479576
rect 45020 479572 45026 479574
rect 117957 479571 118023 479574
rect 147765 479634 147831 479637
rect 213310 479634 213316 479636
rect 147765 479632 213316 479634
rect 147765 479576 147770 479632
rect 147826 479576 213316 479632
rect 147765 479574 213316 479576
rect 147765 479571 147831 479574
rect 213310 479572 213316 479574
rect 213380 479572 213386 479636
rect 233325 479634 233391 479637
rect 364374 479634 364380 479636
rect 233325 479632 364380 479634
rect 233325 479576 233330 479632
rect 233386 479576 364380 479632
rect 233325 479574 364380 479576
rect 233325 479571 233391 479574
rect 364374 479572 364380 479574
rect 364444 479572 364450 479636
rect 44766 479436 44772 479500
rect 44836 479498 44842 479500
rect 118877 479498 118943 479501
rect 44836 479496 118943 479498
rect 44836 479440 118882 479496
rect 118938 479440 118943 479496
rect 44836 479438 118943 479440
rect 44836 479436 44842 479438
rect 118877 479435 118943 479438
rect 154021 479498 154087 479501
rect 208342 479498 208348 479500
rect 154021 479496 208348 479498
rect 154021 479440 154026 479496
rect 154082 479440 208348 479496
rect 154021 479438 208348 479440
rect 154021 479435 154087 479438
rect 208342 479436 208348 479438
rect 208412 479436 208418 479500
rect 210366 479436 210372 479500
rect 210436 479498 210442 479500
rect 512085 479498 512151 479501
rect 210436 479496 512151 479498
rect 210436 479440 512090 479496
rect 512146 479440 512151 479496
rect 210436 479438 512151 479440
rect 210436 479436 210442 479438
rect 512085 479435 512151 479438
rect 152733 478274 152799 478277
rect 209814 478274 209820 478276
rect 152733 478272 209820 478274
rect 152733 478216 152738 478272
rect 152794 478216 209820 478272
rect 152733 478214 209820 478216
rect 152733 478211 152799 478214
rect 209814 478212 209820 478214
rect 209884 478212 209890 478276
rect 223665 478274 223731 478277
rect 378726 478274 378732 478276
rect 223665 478272 378732 478274
rect 223665 478216 223670 478272
rect 223726 478216 378732 478272
rect 223665 478214 378732 478216
rect 223665 478211 223731 478214
rect 378726 478212 378732 478214
rect 378796 478212 378802 478276
rect 62205 478138 62271 478141
rect 198958 478138 198964 478140
rect 62205 478136 198964 478138
rect 62205 478080 62210 478136
rect 62266 478080 198964 478136
rect 62205 478078 198964 478080
rect 62205 478075 62271 478078
rect 198958 478076 198964 478078
rect 199028 478076 199034 478140
rect 204846 478076 204852 478140
rect 204916 478138 204922 478140
rect 457529 478138 457595 478141
rect 204916 478136 457595 478138
rect 204916 478080 457534 478136
rect 457590 478080 457595 478136
rect 204916 478078 457595 478080
rect 204916 478076 204922 478078
rect 457529 478075 457595 478078
rect 43713 477186 43779 477189
rect 124305 477186 124371 477189
rect 43713 477184 124371 477186
rect 43713 477128 43718 477184
rect 43774 477128 124310 477184
rect 124366 477128 124371 477184
rect 43713 477126 124371 477128
rect 43713 477123 43779 477126
rect 124305 477123 124371 477126
rect 43805 477050 43871 477053
rect 125685 477050 125751 477053
rect 43805 477048 125751 477050
rect 43805 476992 43810 477048
rect 43866 476992 125690 477048
rect 125746 476992 125751 477048
rect 43805 476990 125751 476992
rect 43805 476987 43871 476990
rect 125685 476987 125751 476990
rect 297173 477050 297239 477053
rect 376886 477050 376892 477052
rect 297173 477048 376892 477050
rect 297173 476992 297178 477048
rect 297234 476992 376892 477048
rect 297173 476990 376892 476992
rect 297173 476987 297239 476990
rect 376886 476988 376892 476990
rect 376956 476988 376962 477052
rect 43529 476914 43595 476917
rect 125777 476914 125843 476917
rect 43529 476912 125843 476914
rect 43529 476856 43534 476912
rect 43590 476856 125782 476912
rect 125838 476856 125843 476912
rect 43529 476854 125843 476856
rect 43529 476851 43595 476854
rect 125777 476851 125843 476854
rect 145741 476914 145807 476917
rect 203190 476914 203196 476916
rect 145741 476912 203196 476914
rect 145741 476856 145746 476912
rect 145802 476856 203196 476912
rect 145741 476854 203196 476856
rect 145741 476851 145807 476854
rect 203190 476852 203196 476854
rect 203260 476852 203266 476916
rect 227989 476914 228055 476917
rect 370446 476914 370452 476916
rect 227989 476912 370452 476914
rect 227989 476856 227994 476912
rect 228050 476856 370452 476912
rect 227989 476854 370452 476856
rect 227989 476851 228055 476854
rect 370446 476852 370452 476854
rect 370516 476852 370522 476916
rect 43621 476778 43687 476781
rect 127065 476778 127131 476781
rect 43621 476776 127131 476778
rect 43621 476720 43626 476776
rect 43682 476720 127070 476776
rect 127126 476720 127131 476776
rect 43621 476718 127131 476720
rect 43621 476715 43687 476718
rect 127065 476715 127131 476718
rect 151353 476778 151419 476781
rect 214046 476778 214052 476780
rect 151353 476776 214052 476778
rect 151353 476720 151358 476776
rect 151414 476720 214052 476776
rect 151353 476718 214052 476720
rect 151353 476715 151419 476718
rect 214046 476716 214052 476718
rect 214116 476716 214122 476780
rect 234613 476778 234679 476781
rect 378174 476778 378180 476780
rect 234613 476776 378180 476778
rect 234613 476720 234618 476776
rect 234674 476720 378180 476776
rect 234613 476718 378180 476720
rect 234613 476715 234679 476718
rect 378174 476716 378180 476718
rect 378244 476716 378250 476780
rect -960 475540 480 475780
rect 157517 475554 157583 475557
rect 209998 475554 210004 475556
rect 157517 475552 210004 475554
rect 157517 475496 157522 475552
rect 157578 475496 210004 475552
rect 157517 475494 210004 475496
rect 157517 475491 157583 475494
rect 209998 475492 210004 475494
rect 210068 475492 210074 475556
rect 294137 475554 294203 475557
rect 377622 475554 377628 475556
rect 294137 475552 377628 475554
rect 294137 475496 294142 475552
rect 294198 475496 377628 475552
rect 294137 475494 377628 475496
rect 294137 475491 294203 475494
rect 377622 475492 377628 475494
rect 377692 475492 377698 475556
rect 150433 475418 150499 475421
rect 216070 475418 216076 475420
rect 150433 475416 216076 475418
rect 150433 475360 150438 475416
rect 150494 475360 216076 475416
rect 150433 475358 216076 475360
rect 150433 475355 150499 475358
rect 216070 475356 216076 475358
rect 216140 475356 216146 475420
rect 256325 475418 256391 475421
rect 359406 475418 359412 475420
rect 256325 475416 359412 475418
rect 256325 475360 256330 475416
rect 256386 475360 359412 475416
rect 256325 475358 359412 475360
rect 256325 475355 256391 475358
rect 359406 475356 359412 475358
rect 359476 475356 359482 475420
rect 276105 474602 276171 474605
rect 359774 474602 359780 474604
rect 276105 474600 359780 474602
rect 276105 474544 276110 474600
rect 276166 474544 359780 474600
rect 276105 474542 359780 474544
rect 276105 474539 276171 474542
rect 359774 474540 359780 474542
rect 359844 474540 359850 474604
rect 227713 474466 227779 474469
rect 358118 474466 358124 474468
rect 227713 474464 358124 474466
rect 227713 474408 227718 474464
rect 227774 474408 358124 474464
rect 227713 474406 358124 474408
rect 227713 474403 227779 474406
rect 358118 474404 358124 474406
rect 358188 474404 358194 474468
rect 240225 474330 240291 474333
rect 379462 474330 379468 474332
rect 240225 474328 379468 474330
rect 240225 474272 240230 474328
rect 240286 474272 379468 474328
rect 240225 474270 379468 474272
rect 240225 474267 240291 474270
rect 379462 474268 379468 474270
rect 379532 474268 379538 474332
rect 230749 474194 230815 474197
rect 374678 474194 374684 474196
rect 230749 474192 374684 474194
rect 230749 474136 230754 474192
rect 230810 474136 374684 474192
rect 230749 474134 374684 474136
rect 230749 474131 230815 474134
rect 374678 474132 374684 474134
rect 374748 474132 374754 474196
rect 143625 474058 143691 474061
rect 214414 474058 214420 474060
rect 143625 474056 214420 474058
rect 143625 474000 143630 474056
rect 143686 474000 214420 474056
rect 143625 473998 214420 474000
rect 143625 473995 143691 473998
rect 214414 473996 214420 473998
rect 214484 473996 214490 474060
rect 223573 474058 223639 474061
rect 378910 474058 378916 474060
rect 223573 474056 378916 474058
rect 223573 474000 223578 474056
rect 223634 474000 378916 474056
rect 223573 473998 378916 474000
rect 223573 473995 223639 473998
rect 378910 473996 378916 473998
rect 378980 473996 378986 474060
rect 171225 472834 171291 472837
rect 205214 472834 205220 472836
rect 171225 472832 205220 472834
rect 171225 472776 171230 472832
rect 171286 472776 205220 472832
rect 171225 472774 205220 472776
rect 171225 472771 171291 472774
rect 205214 472772 205220 472774
rect 205284 472772 205290 472836
rect 169845 472698 169911 472701
rect 206318 472698 206324 472700
rect 169845 472696 206324 472698
rect 169845 472640 169850 472696
rect 169906 472640 206324 472696
rect 169845 472638 206324 472640
rect 169845 472635 169911 472638
rect 206318 472636 206324 472638
rect 206388 472636 206394 472700
rect 366357 472698 366423 472701
rect 506606 472698 506612 472700
rect 366357 472696 506612 472698
rect 366357 472640 366362 472696
rect 366418 472640 506612 472696
rect 366357 472638 506612 472640
rect 366357 472635 366423 472638
rect 506606 472636 506612 472638
rect 506676 472636 506682 472700
rect 143533 472562 143599 472565
rect 202086 472562 202092 472564
rect 143533 472560 202092 472562
rect 143533 472504 143538 472560
rect 143594 472504 202092 472560
rect 143533 472502 202092 472504
rect 143533 472499 143599 472502
rect 202086 472500 202092 472502
rect 202156 472500 202162 472564
rect 229093 472562 229159 472565
rect 379094 472562 379100 472564
rect 229093 472560 379100 472562
rect 229093 472504 229098 472560
rect 229154 472504 379100 472560
rect 229093 472502 379100 472504
rect 229093 472499 229159 472502
rect 379094 472500 379100 472502
rect 379164 472500 379170 472564
rect 59813 471746 59879 471749
rect 92657 471746 92723 471749
rect 59813 471744 92723 471746
rect 59813 471688 59818 471744
rect 59874 471688 92662 471744
rect 92718 471688 92723 471744
rect 59813 471686 92723 471688
rect 59813 471683 59879 471686
rect 92657 471683 92723 471686
rect 169937 471746 170003 471749
rect 202454 471746 202460 471748
rect 169937 471744 202460 471746
rect 169937 471688 169942 471744
rect 169998 471688 202460 471744
rect 169937 471686 202460 471688
rect 169937 471683 170003 471686
rect 202454 471684 202460 471686
rect 202524 471684 202530 471748
rect 55121 471610 55187 471613
rect 88425 471610 88491 471613
rect 55121 471608 88491 471610
rect 55121 471552 55126 471608
rect 55182 471552 88430 471608
rect 88486 471552 88491 471608
rect 55121 471550 88491 471552
rect 55121 471547 55187 471550
rect 88425 471547 88491 471550
rect 169753 471610 169819 471613
rect 207974 471610 207980 471612
rect 169753 471608 207980 471610
rect 169753 471552 169758 471608
rect 169814 471552 207980 471608
rect 169753 471550 207980 471552
rect 169753 471547 169819 471550
rect 207974 471548 207980 471550
rect 208044 471548 208050 471612
rect 47894 471412 47900 471476
rect 47964 471474 47970 471476
rect 81525 471474 81591 471477
rect 47964 471472 81591 471474
rect 47964 471416 81530 471472
rect 81586 471416 81591 471472
rect 47964 471414 81591 471416
rect 47964 471412 47970 471414
rect 81525 471411 81591 471414
rect 174813 471474 174879 471477
rect 217358 471474 217364 471476
rect 174813 471472 217364 471474
rect 174813 471416 174818 471472
rect 174874 471416 217364 471472
rect 174813 471414 217364 471416
rect 174813 471411 174879 471414
rect 217358 471412 217364 471414
rect 217428 471412 217434 471476
rect 56133 471338 56199 471341
rect 89805 471338 89871 471341
rect 56133 471336 89871 471338
rect 56133 471280 56138 471336
rect 56194 471280 89810 471336
rect 89866 471280 89871 471336
rect 56133 471278 89871 471280
rect 56133 471275 56199 471278
rect 89805 471275 89871 471278
rect 161565 471338 161631 471341
rect 204897 471338 204963 471341
rect 161565 471336 204963 471338
rect 161565 471280 161570 471336
rect 161626 471280 204902 471336
rect 204958 471280 204963 471336
rect 583520 471324 584960 471564
rect 161565 471278 204963 471280
rect 161565 471275 161631 471278
rect 204897 471275 204963 471278
rect 49509 471202 49575 471205
rect 94221 471202 94287 471205
rect 49509 471200 94287 471202
rect 49509 471144 49514 471200
rect 49570 471144 94226 471200
rect 94282 471144 94287 471200
rect 49509 471142 94287 471144
rect 49509 471139 49575 471142
rect 94221 471139 94287 471142
rect 171133 471202 171199 471205
rect 214598 471202 214604 471204
rect 171133 471200 214604 471202
rect 171133 471144 171138 471200
rect 171194 471144 214604 471200
rect 171133 471142 214604 471144
rect 171133 471139 171199 471142
rect 214598 471140 214604 471142
rect 214668 471140 214674 471204
rect 58934 469780 58940 469844
rect 59004 469842 59010 469844
rect 67817 469842 67883 469845
rect 59004 469840 67883 469842
rect 59004 469784 67822 469840
rect 67878 469784 67883 469840
rect 59004 469782 67883 469784
rect 59004 469780 59010 469782
rect 67817 469779 67883 469782
rect 147673 469842 147739 469845
rect 205030 469842 205036 469844
rect 147673 469840 205036 469842
rect 147673 469784 147678 469840
rect 147734 469784 205036 469840
rect 147673 469782 205036 469784
rect 147673 469779 147739 469782
rect 205030 469780 205036 469782
rect 205100 469780 205106 469844
rect 58750 469100 58756 469164
rect 58820 469162 58826 469164
rect 67725 469162 67791 469165
rect 58820 469160 67791 469162
rect 58820 469104 67730 469160
rect 67786 469104 67791 469160
rect 58820 469102 67791 469104
rect 58820 469100 58826 469102
rect 67725 469099 67791 469102
rect 199510 469100 199516 469164
rect 199580 469162 199586 469164
rect 209957 469162 210023 469165
rect 199580 469160 210023 469162
rect 199580 469104 209962 469160
rect 210018 469104 210023 469160
rect 199580 469102 210023 469104
rect 199580 469100 199586 469102
rect 209957 469099 210023 469102
rect 48078 468964 48084 469028
rect 48148 469026 48154 469028
rect 69197 469026 69263 469029
rect 48148 469024 69263 469026
rect 48148 468968 69202 469024
rect 69258 468968 69263 469024
rect 48148 468966 69263 468968
rect 48148 468964 48154 468966
rect 69197 468963 69263 468966
rect 172513 469026 172579 469029
rect 200982 469026 200988 469028
rect 172513 469024 200988 469026
rect 172513 468968 172518 469024
rect 172574 468968 200988 469024
rect 172513 468966 200988 468968
rect 172513 468963 172579 468966
rect 200982 468964 200988 468966
rect 201052 468964 201058 469028
rect 52310 468828 52316 468892
rect 52380 468890 52386 468892
rect 78673 468890 78739 468893
rect 52380 468888 78739 468890
rect 52380 468832 78678 468888
rect 78734 468832 78739 468888
rect 52380 468830 78739 468832
rect 52380 468828 52386 468830
rect 78673 468827 78739 468830
rect 167085 468890 167151 468893
rect 203006 468890 203012 468892
rect 167085 468888 203012 468890
rect 167085 468832 167090 468888
rect 167146 468832 203012 468888
rect 167085 468830 203012 468832
rect 167085 468827 167151 468830
rect 203006 468828 203012 468830
rect 203076 468828 203082 468892
rect 50838 468692 50844 468756
rect 50908 468754 50914 468756
rect 78765 468754 78831 468757
rect 50908 468752 78831 468754
rect 50908 468696 78770 468752
rect 78826 468696 78831 468752
rect 50908 468694 78831 468696
rect 50908 468692 50914 468694
rect 78765 468691 78831 468694
rect 168557 468754 168623 468757
rect 211981 468754 212047 468757
rect 168557 468752 212047 468754
rect 168557 468696 168562 468752
rect 168618 468696 211986 468752
rect 212042 468696 212047 468752
rect 168557 468694 212047 468696
rect 168557 468691 168623 468694
rect 211981 468691 212047 468694
rect 50654 468556 50660 468620
rect 50724 468618 50730 468620
rect 78857 468618 78923 468621
rect 50724 468616 78923 468618
rect 50724 468560 78862 468616
rect 78918 468560 78923 468616
rect 50724 468558 78923 468560
rect 50724 468556 50730 468558
rect 78857 468555 78923 468558
rect 168373 468618 168439 468621
rect 213494 468618 213500 468620
rect 168373 468616 213500 468618
rect 168373 468560 168378 468616
rect 168434 468560 213500 468616
rect 168373 468558 213500 468560
rect 168373 468555 168439 468558
rect 213494 468556 213500 468558
rect 213564 468556 213570 468620
rect 48630 468420 48636 468484
rect 48700 468482 48706 468484
rect 80237 468482 80303 468485
rect 48700 468480 80303 468482
rect 48700 468424 80242 468480
rect 80298 468424 80303 468480
rect 48700 468422 80303 468424
rect 48700 468420 48706 468422
rect 80237 468419 80303 468422
rect 161473 468482 161539 468485
rect 208158 468482 208164 468484
rect 161473 468480 208164 468482
rect 161473 468424 161478 468480
rect 161534 468424 208164 468480
rect 161473 468422 208164 468424
rect 161473 468419 161539 468422
rect 208158 468420 208164 468422
rect 208228 468420 208234 468484
rect 265065 468482 265131 468485
rect 359590 468482 359596 468484
rect 265065 468480 359596 468482
rect 265065 468424 265070 468480
rect 265126 468424 359596 468480
rect 265065 468422 359596 468424
rect 265065 468419 265131 468422
rect 359590 468420 359596 468422
rect 359660 468420 359666 468484
rect 60222 467196 60228 467260
rect 60292 467258 60298 467260
rect 73153 467258 73219 467261
rect 60292 467256 73219 467258
rect 60292 467200 73158 467256
rect 73214 467200 73219 467256
rect 60292 467198 73219 467200
rect 60292 467196 60298 467198
rect 73153 467195 73219 467198
rect 179638 467196 179644 467260
rect 179708 467258 179714 467260
rect 180149 467258 180215 467261
rect 179708 467256 180215 467258
rect 179708 467200 180154 467256
rect 180210 467200 180215 467256
rect 179708 467198 180215 467200
rect 179708 467196 179714 467198
rect 180149 467195 180215 467198
rect 44030 467060 44036 467124
rect 44100 467122 44106 467124
rect 71865 467122 71931 467125
rect 44100 467120 71931 467122
rect 44100 467064 71870 467120
rect 71926 467064 71931 467120
rect 44100 467062 71931 467064
rect 44100 467060 44106 467062
rect 71865 467059 71931 467062
rect 155953 467122 156019 467125
rect 218646 467122 218652 467124
rect 155953 467120 218652 467122
rect 155953 467064 155958 467120
rect 156014 467064 218652 467120
rect 155953 467062 218652 467064
rect 155953 467059 156019 467062
rect 218646 467060 218652 467062
rect 218716 467060 218722 467124
rect 292573 467122 292639 467125
rect 359958 467122 359964 467124
rect 292573 467120 359964 467122
rect 292573 467064 292578 467120
rect 292634 467064 359964 467120
rect 292573 467062 359964 467064
rect 292573 467059 292639 467062
rect 359958 467060 359964 467062
rect 360028 467060 360034 467124
rect 178033 466578 178099 466581
rect 190913 466580 190979 466581
rect 338481 466580 338547 466581
rect 339769 466580 339835 466581
rect 350993 466580 351059 466581
rect 178350 466578 178356 466580
rect 178033 466576 178356 466578
rect 178033 466520 178038 466576
rect 178094 466520 178356 466576
rect 178033 466518 178356 466520
rect 178033 466515 178099 466518
rect 178350 466516 178356 466518
rect 178420 466516 178426 466580
rect 190862 466578 190868 466580
rect 190822 466518 190868 466578
rect 190932 466576 190979 466580
rect 338430 466578 338436 466580
rect 190974 466520 190979 466576
rect 190862 466516 190868 466518
rect 190932 466516 190979 466520
rect 338390 466518 338436 466578
rect 338500 466576 338547 466580
rect 339718 466578 339724 466580
rect 338542 466520 338547 466576
rect 338430 466516 338436 466518
rect 338500 466516 338547 466520
rect 339678 466518 339724 466578
rect 339788 466576 339835 466580
rect 350942 466578 350948 466580
rect 339830 466520 339835 466576
rect 339718 466516 339724 466518
rect 339788 466516 339835 466520
rect 350902 466518 350948 466578
rect 351012 466576 351059 466580
rect 351054 466520 351059 466576
rect 350942 466516 350948 466518
rect 351012 466516 351059 466520
rect 190913 466515 190979 466516
rect 338481 466515 338547 466516
rect 339769 466515 339835 466516
rect 350993 466515 351059 466516
rect 498469 466580 498535 466581
rect 499757 466580 499823 466581
rect 510889 466580 510955 466581
rect 498469 466576 498516 466580
rect 498580 466578 498586 466580
rect 498469 466520 498474 466576
rect 498469 466516 498516 466520
rect 498580 466518 498626 466578
rect 499757 466576 499804 466580
rect 499868 466578 499874 466580
rect 510838 466578 510844 466580
rect 499757 466520 499762 466576
rect 498580 466516 498586 466518
rect 499757 466516 499804 466520
rect 499868 466518 499914 466578
rect 510798 466518 510844 466578
rect 510908 466576 510955 466580
rect 510950 466520 510955 466576
rect 499868 466516 499874 466518
rect 510838 466516 510844 466518
rect 510908 466516 510955 466520
rect 498469 466515 498535 466516
rect 499757 466515 499823 466516
rect 510889 466515 510955 466516
rect 50470 466380 50476 466444
rect 50540 466442 50546 466444
rect 66253 466442 66319 466445
rect 50540 466440 66319 466442
rect 50540 466384 66258 466440
rect 66314 466384 66319 466440
rect 50540 466382 66319 466384
rect 50540 466380 50546 466382
rect 66253 466379 66319 466382
rect 55070 466244 55076 466308
rect 55140 466306 55146 466308
rect 71773 466306 71839 466309
rect 55140 466304 71839 466306
rect 55140 466248 71778 466304
rect 71834 466248 71839 466304
rect 55140 466246 71839 466248
rect 55140 466244 55146 466246
rect 71773 466243 71839 466246
rect 182817 466306 182883 466309
rect 198774 466306 198780 466308
rect 182817 466304 198780 466306
rect 182817 466248 182822 466304
rect 182878 466248 198780 466304
rect 182817 466246 198780 466248
rect 182817 466243 182883 466246
rect 198774 466244 198780 466246
rect 198844 466244 198850 466308
rect 55438 466108 55444 466172
rect 55508 466170 55514 466172
rect 74533 466170 74599 466173
rect 55508 466168 74599 466170
rect 55508 466112 74538 466168
rect 74594 466112 74599 466168
rect 55508 466110 74599 466112
rect 55508 466108 55514 466110
rect 74533 466107 74599 466110
rect 165797 466170 165863 466173
rect 204989 466170 205055 466173
rect 165797 466168 205055 466170
rect 165797 466112 165802 466168
rect 165858 466112 204994 466168
rect 205050 466112 205055 466168
rect 165797 466110 205055 466112
rect 165797 466107 165863 466110
rect 204989 466107 205055 466110
rect 54886 465972 54892 466036
rect 54956 466034 54962 466036
rect 76005 466034 76071 466037
rect 54956 466032 76071 466034
rect 54956 465976 76010 466032
rect 76066 465976 76071 466032
rect 54956 465974 76071 465976
rect 54956 465972 54962 465974
rect 76005 465971 76071 465974
rect 166993 466034 167059 466037
rect 206461 466034 206527 466037
rect 166993 466032 206527 466034
rect 166993 465976 166998 466032
rect 167054 465976 206466 466032
rect 206522 465976 206527 466032
rect 166993 465974 206527 465976
rect 166993 465971 167059 465974
rect 206461 465971 206527 465974
rect 46606 465836 46612 465900
rect 46676 465898 46682 465900
rect 69013 465898 69079 465901
rect 46676 465896 69079 465898
rect 46676 465840 69018 465896
rect 69074 465840 69079 465896
rect 46676 465838 69079 465840
rect 46676 465836 46682 465838
rect 69013 465835 69079 465838
rect 162853 465898 162919 465901
rect 216121 465898 216187 465901
rect 162853 465896 216187 465898
rect 162853 465840 162858 465896
rect 162914 465840 216126 465896
rect 216182 465840 216187 465896
rect 162853 465838 216187 465840
rect 162853 465835 162919 465838
rect 216121 465835 216187 465838
rect 52126 465700 52132 465764
rect 52196 465762 52202 465764
rect 74625 465762 74691 465765
rect 52196 465760 74691 465762
rect 52196 465704 74630 465760
rect 74686 465704 74691 465760
rect 52196 465702 74691 465704
rect 52196 465700 52202 465702
rect 74625 465699 74691 465702
rect 165613 465762 165679 465765
rect 218973 465762 219039 465765
rect 165613 465760 219039 465762
rect 165613 465704 165618 465760
rect 165674 465704 218978 465760
rect 219034 465704 219039 465760
rect 165613 465702 219039 465704
rect 165613 465699 165679 465702
rect 218973 465699 219039 465702
rect 58566 465564 58572 465628
rect 58636 465626 58642 465628
rect 69105 465626 69171 465629
rect 58636 465624 69171 465626
rect 58636 465568 69110 465624
rect 69166 465568 69171 465624
rect 58636 465566 69171 465568
rect 58636 465564 58642 465566
rect 69105 465563 69171 465566
rect 51574 465156 51580 465220
rect 51644 465218 51650 465220
rect 51993 465218 52059 465221
rect 55673 465220 55739 465221
rect 55622 465218 55628 465220
rect 51644 465216 52059 465218
rect 51644 465160 51998 465216
rect 52054 465160 52059 465216
rect 51644 465158 52059 465160
rect 55582 465158 55628 465218
rect 55692 465216 55739 465220
rect 55734 465160 55739 465216
rect 51644 465156 51650 465158
rect 51993 465155 52059 465158
rect 55622 465156 55628 465158
rect 55692 465156 55739 465160
rect 55673 465155 55739 465156
rect 125593 464402 125659 464405
rect 199142 464402 199148 464404
rect 125593 464400 199148 464402
rect 125593 464344 125598 464400
rect 125654 464344 199148 464400
rect 125593 464342 199148 464344
rect 125593 464339 125659 464342
rect 199142 464340 199148 464342
rect 199212 464340 199218 464404
rect -960 462634 480 462724
rect 3693 462634 3759 462637
rect -960 462632 3759 462634
rect -960 462576 3698 462632
rect 3754 462576 3759 462632
rect -960 462574 3759 462576
rect -960 462484 480 462574
rect 3693 462571 3759 462574
rect 196558 460186 196618 460190
rect 198917 460186 198983 460189
rect 196558 460184 198983 460186
rect 196558 460128 198922 460184
rect 198978 460128 198983 460184
rect 196558 460126 198983 460128
rect 356562 460186 356622 460190
rect 358813 460186 358879 460189
rect 356562 460184 358879 460186
rect 356562 460128 358818 460184
rect 358874 460128 358879 460184
rect 356562 460126 358879 460128
rect 198917 460123 198983 460126
rect 358813 460123 358879 460126
rect 516558 459642 516618 460190
rect 518893 459642 518959 459645
rect 519445 459642 519511 459645
rect 516558 459640 519511 459642
rect 516558 459584 518898 459640
rect 518954 459584 519450 459640
rect 519506 459584 519511 459640
rect 516558 459582 519511 459584
rect 518893 459579 518959 459582
rect 519445 459579 519511 459582
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect 57881 417346 57947 417349
rect 60002 417346 60062 417894
rect 216673 417890 216739 417893
rect 219390 417890 220064 417924
rect 216673 417888 220064 417890
rect 216673 417832 216678 417888
rect 216734 417864 220064 417888
rect 376937 417890 377003 417893
rect 379470 417890 380052 417924
rect 376937 417888 380052 417890
rect 216734 417832 219450 417864
rect 216673 417830 219450 417832
rect 376937 417832 376942 417888
rect 376998 417864 380052 417888
rect 376998 417832 379530 417864
rect 376937 417830 379530 417832
rect 216673 417827 216739 417830
rect 376937 417827 377003 417830
rect 57881 417344 60062 417346
rect 57881 417288 57886 417344
rect 57942 417288 60062 417344
rect 57881 417286 60062 417288
rect 57881 417283 57947 417286
rect 56961 417210 57027 417213
rect 56961 417208 60062 417210
rect 56961 417152 56966 417208
rect 57022 417152 60062 417208
rect 56961 417150 60062 417152
rect 56961 417147 57027 417150
rect 60002 416942 60062 417150
rect 217961 416938 218027 416941
rect 219390 416938 220064 416972
rect 217961 416936 220064 416938
rect 217961 416880 217966 416936
rect 218022 416912 220064 416936
rect 377765 416938 377831 416941
rect 379470 416938 380052 416972
rect 377765 416936 380052 416938
rect 218022 416880 219450 416912
rect 217961 416878 219450 416880
rect 377765 416880 377770 416936
rect 377826 416912 380052 416936
rect 377826 416880 379530 416912
rect 377765 416878 379530 416880
rect 217961 416875 218027 416878
rect 377765 416875 377831 416878
rect 57881 414218 57947 414221
rect 60002 414218 60062 414766
rect 217133 414762 217199 414765
rect 219390 414762 220064 414796
rect 217133 414760 220064 414762
rect 217133 414704 217138 414760
rect 217194 414736 220064 414760
rect 377673 414762 377739 414765
rect 379470 414762 380052 414796
rect 377673 414760 380052 414762
rect 217194 414704 219450 414736
rect 217133 414702 219450 414704
rect 377673 414704 377678 414760
rect 377734 414736 380052 414760
rect 377734 414704 379530 414736
rect 377673 414702 379530 414704
rect 217133 414699 217199 414702
rect 377673 414699 377739 414702
rect 57881 414216 60062 414218
rect 57881 414160 57886 414216
rect 57942 414160 60062 414216
rect 57881 414158 60062 414160
rect 57881 414155 57947 414158
rect 57881 413266 57947 413269
rect 60002 413266 60062 413814
rect 216857 413810 216923 413813
rect 219390 413810 220064 413844
rect 216857 413808 220064 413810
rect 216857 413752 216862 413808
rect 216918 413784 220064 413808
rect 377765 413810 377831 413813
rect 379470 413810 380052 413844
rect 377765 413808 380052 413810
rect 216918 413752 219450 413784
rect 216857 413750 219450 413752
rect 377765 413752 377770 413808
rect 377826 413784 380052 413808
rect 377826 413752 379530 413784
rect 377765 413750 379530 413752
rect 216857 413747 216923 413750
rect 377765 413747 377831 413750
rect 57881 413264 60062 413266
rect 57881 413208 57886 413264
rect 57942 413208 60062 413264
rect 57881 413206 60062 413208
rect 57881 413203 57947 413206
rect 57881 411498 57947 411501
rect 60002 411498 60062 412046
rect 217685 412042 217751 412045
rect 219390 412042 220064 412076
rect 217685 412040 220064 412042
rect 217685 411984 217690 412040
rect 217746 412016 220064 412040
rect 377029 412042 377095 412045
rect 377581 412042 377647 412045
rect 379470 412042 380052 412076
rect 377029 412040 380052 412042
rect 217746 411984 219450 412016
rect 217685 411982 219450 411984
rect 377029 411984 377034 412040
rect 377090 411984 377586 412040
rect 377642 412016 380052 412040
rect 377642 411984 379530 412016
rect 377029 411982 379530 411984
rect 217685 411979 217751 411982
rect 377029 411979 377095 411982
rect 377581 411979 377647 411982
rect 57881 411496 60062 411498
rect 57881 411440 57886 411496
rect 57942 411440 60062 411496
rect 57881 411438 60062 411440
rect 57881 411435 57947 411438
rect 205398 411300 205404 411364
rect 205468 411362 205474 411364
rect 205541 411362 205607 411365
rect 205468 411360 205607 411362
rect 205468 411304 205546 411360
rect 205602 411304 205607 411360
rect 205468 411302 205607 411304
rect 205468 411300 205474 411302
rect 205541 411299 205607 411302
rect 217225 411362 217291 411365
rect 217685 411362 217751 411365
rect 217225 411360 217751 411362
rect 217225 411304 217230 411360
rect 217286 411304 217690 411360
rect 217746 411304 217751 411360
rect 217225 411302 217751 411304
rect 217225 411299 217291 411302
rect 217685 411299 217751 411302
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 57881 410410 57947 410413
rect 60002 410410 60062 410958
rect 216765 410954 216831 410957
rect 219390 410954 220064 410988
rect 216765 410952 220064 410954
rect 216765 410896 216770 410952
rect 216826 410928 220064 410952
rect 377029 410954 377095 410957
rect 379470 410954 380052 410988
rect 377029 410952 380052 410954
rect 216826 410896 219450 410928
rect 216765 410894 219450 410896
rect 377029 410896 377034 410952
rect 377090 410928 380052 410952
rect 377090 410896 379530 410928
rect 377029 410894 379530 410896
rect 216765 410891 216831 410894
rect 377029 410891 377095 410894
rect 57881 410408 60062 410410
rect 57881 410352 57886 410408
rect 57942 410352 60062 410408
rect 57881 410350 60062 410352
rect 57881 410347 57947 410350
rect 57881 408642 57947 408645
rect 60002 408642 60062 409190
rect 217317 409186 217383 409189
rect 217869 409186 217935 409189
rect 219390 409186 220064 409220
rect 217317 409184 220064 409186
rect 217317 409128 217322 409184
rect 217378 409128 217874 409184
rect 217930 409160 220064 409184
rect 377397 409186 377463 409189
rect 378041 409186 378107 409189
rect 379470 409186 380052 409220
rect 377397 409184 380052 409186
rect 217930 409128 219450 409160
rect 217317 409126 219450 409128
rect 377397 409128 377402 409184
rect 377458 409128 378046 409184
rect 378102 409160 380052 409184
rect 378102 409128 379530 409160
rect 377397 409126 379530 409128
rect 217317 409123 217383 409126
rect 217869 409123 217935 409126
rect 377397 409123 377463 409126
rect 378041 409123 378107 409126
rect 57881 408640 60062 408642
rect 57881 408584 57886 408640
rect 57942 408584 60062 408640
rect 57881 408582 60062 408584
rect 57881 408579 57947 408582
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 196558 400346 196618 400350
rect 199561 400346 199627 400349
rect 196558 400344 199627 400346
rect 196558 400288 199566 400344
rect 199622 400288 199627 400344
rect 196558 400286 199627 400288
rect 356562 400346 356622 400350
rect 358905 400346 358971 400349
rect 356562 400344 358971 400346
rect 356562 400288 358910 400344
rect 358966 400288 358971 400344
rect 356562 400286 358971 400288
rect 516558 400346 516618 400350
rect 519077 400346 519143 400349
rect 516558 400344 519143 400346
rect 516558 400288 519082 400344
rect 519138 400288 519143 400344
rect 516558 400286 519143 400288
rect 199561 400283 199627 400286
rect 358905 400283 358971 400286
rect 519077 400283 519143 400286
rect 196558 398170 196618 398718
rect 199193 398170 199259 398173
rect 196558 398168 199259 398170
rect 196558 398112 199198 398168
rect 199254 398112 199259 398168
rect 196558 398110 199259 398112
rect 356562 398170 356622 398718
rect 358997 398170 359063 398173
rect 356562 398168 359063 398170
rect 356562 398112 359002 398168
rect 359058 398112 359063 398168
rect 356562 398110 359063 398112
rect 516558 398170 516618 398718
rect 518985 398170 519051 398173
rect 516558 398168 519051 398170
rect 516558 398112 518990 398168
rect 519046 398112 519051 398168
rect 516558 398110 519051 398112
rect 199193 398107 199259 398110
rect 358997 398107 359063 398110
rect 518985 398107 519051 398110
rect 198181 398034 198247 398037
rect 199142 398034 199148 398036
rect 198181 398032 199148 398034
rect 198181 397976 198186 398032
rect 198242 397976 199148 398032
rect 198181 397974 199148 397976
rect 198181 397971 198247 397974
rect 199142 397972 199148 397974
rect 199212 397972 199218 398036
rect -960 397340 480 397580
rect 196558 396810 196618 397358
rect 199101 396810 199167 396813
rect 196558 396808 199167 396810
rect 196558 396752 199106 396808
rect 199162 396752 199167 396808
rect 196558 396750 199167 396752
rect 356562 396810 356622 397358
rect 359825 396810 359891 396813
rect 356562 396808 359891 396810
rect 356562 396752 359830 396808
rect 359886 396752 359891 396808
rect 356562 396750 359891 396752
rect 516558 396810 516618 397358
rect 519169 396810 519235 396813
rect 516558 396808 519235 396810
rect 516558 396752 519174 396808
rect 519230 396752 519235 396808
rect 516558 396750 519235 396752
rect 199101 396747 199167 396750
rect 359825 396747 359891 396750
rect 519169 396747 519235 396750
rect 199193 396132 199259 396133
rect 199142 396130 199148 396132
rect 199102 396070 199148 396130
rect 199212 396128 199259 396132
rect 199254 396072 199259 396128
rect 199142 396068 199148 396070
rect 199212 396068 199259 396072
rect 199193 396067 199259 396068
rect 196558 395858 196618 395862
rect 199326 395858 199332 395860
rect 196558 395798 199332 395858
rect 199326 395796 199332 395798
rect 199396 395796 199402 395860
rect 356562 395314 356622 395862
rect 359917 395314 359983 395317
rect 356562 395312 359983 395314
rect 356562 395256 359922 395312
rect 359978 395256 359983 395312
rect 356562 395254 359983 395256
rect 516558 395314 516618 395862
rect 519353 395314 519419 395317
rect 516558 395312 519419 395314
rect 516558 395256 519358 395312
rect 519414 395256 519419 395312
rect 516558 395254 519419 395256
rect 359917 395251 359983 395254
rect 519353 395251 519419 395254
rect 196558 394634 196618 394638
rect 199745 394634 199811 394637
rect 196558 394632 199811 394634
rect 196558 394576 199750 394632
rect 199806 394576 199811 394632
rect 196558 394574 199811 394576
rect 199745 394571 199811 394574
rect 356562 394090 356622 394638
rect 359089 394090 359155 394093
rect 356562 394088 359155 394090
rect 356562 394032 359094 394088
rect 359150 394032 359155 394088
rect 356562 394030 359155 394032
rect 516558 394090 516618 394638
rect 519261 394090 519327 394093
rect 516558 394088 519327 394090
rect 516558 394032 519266 394088
rect 519322 394032 519327 394088
rect 516558 394030 519327 394032
rect 359089 394027 359155 394030
rect 519261 394027 519327 394030
rect 583520 391628 584960 391868
rect 57053 391506 57119 391509
rect 57053 391504 60062 391506
rect 57053 391448 57058 391504
rect 57114 391448 60062 391504
rect 57053 391446 60062 391448
rect 57053 391443 57119 391446
rect 60002 390966 60062 391446
rect 216673 390962 216739 390965
rect 219390 390962 220064 390996
rect 216673 390960 220064 390962
rect 216673 390904 216678 390960
rect 216734 390936 220064 390960
rect 376937 390962 377003 390965
rect 379470 390962 380052 390996
rect 376937 390960 380052 390962
rect 216734 390904 219450 390936
rect 216673 390902 219450 390904
rect 376937 390904 376942 390960
rect 376998 390936 380052 390960
rect 376998 390904 379530 390936
rect 376937 390902 379530 390904
rect 216673 390899 216739 390902
rect 376937 390899 377003 390902
rect 208342 390628 208348 390692
rect 208412 390690 208418 390692
rect 208669 390690 208735 390693
rect 208412 390688 208735 390690
rect 208412 390632 208674 390688
rect 208730 390632 208735 390688
rect 208412 390630 208735 390632
rect 208412 390628 208418 390630
rect 208669 390627 208735 390630
rect 57513 389330 57579 389333
rect 59494 389330 60032 389364
rect 57513 389328 60032 389330
rect 57513 389272 57518 389328
rect 57574 389304 60032 389328
rect 216673 389330 216739 389333
rect 219390 389330 220064 389364
rect 216673 389328 220064 389330
rect 57574 389272 59554 389304
rect 57513 389270 59554 389272
rect 216673 389272 216678 389328
rect 216734 389304 220064 389328
rect 376937 389330 377003 389333
rect 379470 389330 380052 389364
rect 376937 389328 380052 389330
rect 216734 389272 219450 389304
rect 216673 389270 219450 389272
rect 376937 389272 376942 389328
rect 376998 389304 380052 389328
rect 376998 389272 379530 389304
rect 376937 389270 379530 389272
rect 57513 389267 57579 389270
rect 216673 389267 216739 389270
rect 376937 389267 377003 389270
rect 57053 389058 57119 389061
rect 60002 389058 60062 389062
rect 57053 389056 60062 389058
rect 57053 389000 57058 389056
rect 57114 389000 60062 389056
rect 57053 388998 60062 389000
rect 216673 389058 216739 389061
rect 219390 389058 220064 389092
rect 216673 389056 220064 389058
rect 216673 389000 216678 389056
rect 216734 389032 220064 389056
rect 376937 389058 377003 389061
rect 379470 389058 380052 389092
rect 376937 389056 380052 389058
rect 216734 389000 219450 389032
rect 216673 388998 219450 389000
rect 376937 389000 376942 389056
rect 376998 389032 380052 389056
rect 376998 389000 379530 389032
rect 376937 388998 379530 389000
rect 57053 388995 57119 388998
rect 216673 388995 216739 388998
rect 376937 388995 377003 388998
rect 51942 388452 51948 388516
rect 52012 388514 52018 388516
rect 52361 388514 52427 388517
rect 52012 388512 52427 388514
rect 52012 388456 52366 388512
rect 52422 388456 52427 388512
rect 52012 388454 52427 388456
rect 52012 388452 52018 388454
rect 52361 388451 52427 388454
rect 57646 388452 57652 388516
rect 57716 388514 57722 388516
rect 58617 388514 58683 388517
rect 57716 388512 58683 388514
rect 57716 388456 58622 388512
rect 58678 388456 58683 388512
rect 57716 388454 58683 388456
rect 57716 388452 57722 388454
rect 58617 388451 58683 388454
rect -960 384284 480 384524
rect 377622 382332 377628 382396
rect 377692 382394 377698 382396
rect 379605 382394 379671 382397
rect 377692 382392 379671 382394
rect 377692 382336 379610 382392
rect 379666 382336 379671 382392
rect 377692 382334 379671 382336
rect 377692 382332 377698 382334
rect 379605 382331 379671 382334
rect 359958 381516 359964 381580
rect 360028 381578 360034 381580
rect 374269 381578 374335 381581
rect 375189 381578 375255 381581
rect 360028 381576 375255 381578
rect 360028 381520 374274 381576
rect 374330 381520 375194 381576
rect 375250 381520 375255 381576
rect 360028 381518 375255 381520
rect 360028 381516 360034 381518
rect 374269 381515 374335 381518
rect 375189 381515 375255 381518
rect 59854 380972 59860 381036
rect 59924 381034 59930 381036
rect 59997 381034 60063 381037
rect 59924 381032 60063 381034
rect 59924 380976 60002 381032
rect 60058 380976 60063 381032
rect 59924 380974 60063 380976
rect 59924 380972 59930 380974
rect 59997 380971 60063 380974
rect 205582 380972 205588 381036
rect 205652 381034 205658 381036
rect 206185 381034 206251 381037
rect 205652 381032 206251 381034
rect 205652 380976 206190 381032
rect 206246 380976 206251 381032
rect 205652 380974 206251 380976
rect 205652 380972 205658 380974
rect 206185 380971 206251 380974
rect 93393 380900 93459 380901
rect 110965 380900 111031 380901
rect 113541 380900 113607 380901
rect 116025 380900 116091 380901
rect 118417 380900 118483 380901
rect 120993 380900 121059 380901
rect 93393 380896 93462 380900
rect 93393 380840 93398 380896
rect 93454 380840 93462 380896
rect 93393 380836 93462 380840
rect 93526 380898 93532 380900
rect 93526 380838 93550 380898
rect 110965 380896 111006 380900
rect 111070 380898 111076 380900
rect 110965 380840 110970 380896
rect 93526 380836 93532 380838
rect 110965 380836 111006 380840
rect 111070 380838 111122 380898
rect 113541 380896 113590 380900
rect 113654 380898 113660 380900
rect 113541 380840 113546 380896
rect 111070 380836 111076 380838
rect 113541 380836 113590 380840
rect 113654 380838 113698 380898
rect 116025 380896 116038 380900
rect 116102 380898 116108 380900
rect 116025 380840 116030 380896
rect 113654 380836 113660 380838
rect 116025 380836 116038 380840
rect 116102 380838 116182 380898
rect 118417 380896 118486 380900
rect 118417 380840 118422 380896
rect 118478 380840 118486 380896
rect 116102 380836 116108 380838
rect 118417 380836 118486 380840
rect 118550 380898 118556 380900
rect 120928 380898 120934 380900
rect 118550 380838 118574 380898
rect 120902 380838 120934 380898
rect 118550 380836 118556 380838
rect 120928 380836 120934 380838
rect 120998 380896 121059 380900
rect 121054 380840 121059 380896
rect 120998 380836 121059 380840
rect 93393 380835 93459 380836
rect 110965 380835 111031 380836
rect 113541 380835 113607 380836
rect 116025 380835 116091 380836
rect 118417 380835 118483 380836
rect 120993 380835 121059 380836
rect 123477 380900 123543 380901
rect 125961 380900 126027 380901
rect 131021 380900 131087 380901
rect 133505 380900 133571 380901
rect 135897 380900 135963 380901
rect 143533 380900 143599 380901
rect 146017 380900 146083 380901
rect 158529 380900 158595 380901
rect 160921 380900 160987 380901
rect 163405 380900 163471 380901
rect 165981 380900 166047 380901
rect 123477 380896 123518 380900
rect 123582 380898 123588 380900
rect 123477 380840 123482 380896
rect 123477 380836 123518 380840
rect 123582 380838 123634 380898
rect 123582 380836 123588 380838
rect 125960 380836 125966 380900
rect 126030 380898 126036 380900
rect 130992 380898 130998 380900
rect 126030 380838 126118 380898
rect 130930 380838 130998 380898
rect 131062 380896 131087 380900
rect 133440 380898 133446 380900
rect 131082 380840 131087 380896
rect 126030 380836 126036 380838
rect 130992 380836 130998 380838
rect 131062 380836 131087 380840
rect 133414 380838 133446 380898
rect 133440 380836 133446 380838
rect 133510 380896 133571 380900
rect 135888 380898 135894 380900
rect 133566 380840 133571 380896
rect 133510 380836 133571 380840
rect 135806 380838 135894 380898
rect 135888 380836 135894 380838
rect 135958 380836 135964 380900
rect 143504 380898 143510 380900
rect 143442 380838 143510 380898
rect 143574 380896 143599 380900
rect 145952 380898 145958 380900
rect 143594 380840 143599 380896
rect 143504 380836 143510 380838
rect 143574 380836 143599 380840
rect 145926 380838 145958 380898
rect 145952 380836 145958 380838
rect 146022 380896 146083 380900
rect 158464 380898 158470 380900
rect 146078 380840 146083 380896
rect 146022 380836 146083 380840
rect 158438 380838 158470 380898
rect 158464 380836 158470 380838
rect 158534 380896 158595 380900
rect 160912 380898 160918 380900
rect 158590 380840 158595 380896
rect 158534 380836 158595 380840
rect 160830 380838 160918 380898
rect 160912 380836 160918 380838
rect 160982 380836 160988 380900
rect 163360 380898 163366 380900
rect 163314 380838 163366 380898
rect 163430 380896 163471 380900
rect 165944 380898 165950 380900
rect 163466 380840 163471 380896
rect 163360 380836 163366 380838
rect 163430 380836 163471 380840
rect 165890 380838 165950 380898
rect 166014 380896 166047 380900
rect 166042 380840 166047 380896
rect 165944 380836 165950 380838
rect 166014 380836 166047 380840
rect 123477 380835 123543 380836
rect 125961 380835 126027 380836
rect 131021 380835 131087 380836
rect 133505 380835 133571 380836
rect 135897 380835 135963 380836
rect 143533 380835 143599 380836
rect 146017 380835 146083 380836
rect 158529 380835 158595 380836
rect 160921 380835 160987 380836
rect 163405 380835 163471 380836
rect 165981 380835 166047 380836
rect 215477 380898 215543 380901
rect 216581 380898 216647 380901
rect 263928 380898 263934 380900
rect 215477 380896 263934 380898
rect 215477 380840 215482 380896
rect 215538 380840 216586 380896
rect 216642 380840 263934 380896
rect 215477 380838 263934 380840
rect 215477 380835 215543 380838
rect 216581 380835 216647 380838
rect 263928 380836 263934 380838
rect 263998 380836 264004 380900
rect 376385 380898 376451 380901
rect 485944 380898 485950 380900
rect 376385 380896 485950 380898
rect 376385 380840 376390 380896
rect 376446 380840 485950 380896
rect 376385 380838 485950 380840
rect 376385 380835 376451 380838
rect 485944 380836 485950 380838
rect 486014 380836 486020 380900
rect 50981 380762 51047 380765
rect 216673 380762 216739 380765
rect 50981 380760 216739 380762
rect 50981 380704 50986 380760
rect 51042 380704 216678 380760
rect 216734 380704 216739 380760
rect 50981 380702 216739 380704
rect 50981 380699 51047 380702
rect 216673 380699 216739 380702
rect 235993 380764 236059 380765
rect 237097 380764 237163 380765
rect 243077 380764 243143 380765
rect 245377 380764 245443 380765
rect 256049 380764 256115 380765
rect 269757 380764 269823 380765
rect 421097 380764 421163 380765
rect 422845 380764 422911 380765
rect 430941 380764 431007 380765
rect 433609 380764 433675 380765
rect 235993 380760 236054 380764
rect 235993 380704 235998 380760
rect 235993 380700 236054 380704
rect 236118 380762 236124 380764
rect 236118 380702 236150 380762
rect 237097 380760 237142 380764
rect 237206 380762 237212 380764
rect 237097 380704 237102 380760
rect 236118 380700 236124 380702
rect 237097 380700 237142 380704
rect 237206 380702 237254 380762
rect 243077 380760 243126 380764
rect 243190 380762 243196 380764
rect 243077 380704 243082 380760
rect 237206 380700 237212 380702
rect 243077 380700 243126 380704
rect 243190 380702 243234 380762
rect 245377 380760 245438 380764
rect 245377 380704 245382 380760
rect 243190 380700 243196 380702
rect 245377 380700 245438 380704
rect 245502 380762 245508 380764
rect 256040 380762 256046 380764
rect 245502 380702 245534 380762
rect 255958 380702 256046 380762
rect 245502 380700 245508 380702
rect 256040 380700 256046 380702
rect 256110 380700 256116 380764
rect 269757 380760 269782 380764
rect 269846 380762 269852 380764
rect 421072 380762 421078 380764
rect 269757 380704 269762 380760
rect 269757 380700 269782 380704
rect 269846 380702 269914 380762
rect 421006 380702 421078 380762
rect 421142 380760 421163 380764
rect 422840 380762 422846 380764
rect 421158 380704 421163 380760
rect 269846 380700 269852 380702
rect 421072 380700 421078 380702
rect 421142 380700 421163 380704
rect 422754 380702 422846 380762
rect 422840 380700 422846 380702
rect 422910 380700 422916 380764
rect 430941 380760 431006 380764
rect 430941 380704 430946 380760
rect 431002 380704 431006 380760
rect 430941 380700 431006 380704
rect 431070 380762 431076 380764
rect 433584 380762 433590 380764
rect 431070 380702 431098 380762
rect 433518 380702 433590 380762
rect 433654 380760 433675 380764
rect 433670 380704 433675 380760
rect 431070 380700 431076 380702
rect 433584 380700 433590 380702
rect 433654 380700 433675 380704
rect 235993 380699 236059 380700
rect 237097 380699 237163 380700
rect 243077 380699 243143 380700
rect 245377 380699 245443 380700
rect 256049 380699 256115 380700
rect 269757 380699 269823 380700
rect 421097 380699 421163 380700
rect 422845 380699 422911 380700
rect 430941 380699 431007 380700
rect 433609 380699 433675 380700
rect 436001 380764 436067 380765
rect 438485 380764 438551 380765
rect 440877 380764 440943 380765
rect 443453 380764 443519 380765
rect 436001 380760 436038 380764
rect 436102 380762 436108 380764
rect 438480 380762 438486 380764
rect 436001 380704 436006 380760
rect 436001 380700 436038 380704
rect 436102 380702 436158 380762
rect 438394 380702 438486 380762
rect 436102 380700 436108 380702
rect 438480 380700 438486 380702
rect 438550 380700 438556 380764
rect 440877 380760 440934 380764
rect 440998 380762 441004 380764
rect 440877 380704 440882 380760
rect 440877 380700 440934 380704
rect 440998 380702 441034 380762
rect 443453 380760 443518 380764
rect 443453 380704 443458 380760
rect 443514 380704 443518 380760
rect 440998 380700 441004 380702
rect 443453 380700 443518 380704
rect 443582 380762 443588 380764
rect 443582 380702 443610 380762
rect 443582 380700 443588 380702
rect 436001 380699 436067 380700
rect 438485 380699 438551 380700
rect 440877 380699 440943 380700
rect 443453 380699 443519 380700
rect 77136 380564 77142 380628
rect 77206 380626 77212 380628
rect 204345 380626 204411 380629
rect 254485 380628 254551 380629
rect 255865 380628 255931 380629
rect 256969 380628 257035 380629
rect 259453 380628 259519 380629
rect 265249 380628 265315 380629
rect 270953 380628 271019 380629
rect 408677 380628 408743 380629
rect 413461 380628 413527 380629
rect 419441 380628 419507 380629
rect 434345 380628 434411 380629
rect 445937 380628 446003 380629
rect 77206 380624 204411 380626
rect 77206 380568 204350 380624
rect 204406 380568 204411 380624
rect 77206 380566 204411 380568
rect 77206 380564 77212 380566
rect 204345 380563 204411 380566
rect 219390 380566 253950 380626
rect 76046 380428 76052 380492
rect 76116 380490 76122 380492
rect 76116 380430 200130 380490
rect 76116 380428 76122 380430
rect 128353 380356 128419 380357
rect 155953 380356 156019 380357
rect 128302 380354 128308 380356
rect 128262 380294 128308 380354
rect 128372 380352 128419 380356
rect 155902 380354 155908 380356
rect 128414 380296 128419 380352
rect 128302 380292 128308 380294
rect 128372 380292 128419 380296
rect 155862 380294 155908 380354
rect 155972 380352 156019 380356
rect 156014 380296 156019 380352
rect 155902 380292 155908 380294
rect 155972 380292 156019 380296
rect 200070 380354 200130 380430
rect 216622 380428 216628 380492
rect 216692 380490 216698 380492
rect 216990 380490 216996 380492
rect 216692 380430 216996 380490
rect 216692 380428 216698 380430
rect 216990 380428 216996 380430
rect 217060 380490 217066 380492
rect 219390 380490 219450 380566
rect 217060 380430 219450 380490
rect 253890 380490 253950 380566
rect 254485 380624 254550 380628
rect 254485 380568 254490 380624
rect 254546 380568 254550 380624
rect 254485 380564 254550 380568
rect 254614 380626 254620 380628
rect 254614 380566 254642 380626
rect 255865 380624 255910 380628
rect 255974 380626 255980 380628
rect 255865 380568 255870 380624
rect 254614 380564 254620 380566
rect 255865 380564 255910 380568
rect 255974 380566 256022 380626
rect 256969 380624 256998 380628
rect 257062 380626 257068 380628
rect 259440 380626 259446 380628
rect 256969 380568 256974 380624
rect 255974 380564 255980 380566
rect 256969 380564 256998 380568
rect 257062 380566 257126 380626
rect 259362 380566 259446 380626
rect 259510 380624 259519 380628
rect 259514 380568 259519 380624
rect 257062 380564 257068 380566
rect 259440 380564 259446 380566
rect 259510 380564 259519 380568
rect 260664 380564 260670 380628
rect 260734 380564 260740 380628
rect 265249 380624 265294 380628
rect 265358 380626 265364 380628
rect 265249 380568 265254 380624
rect 265249 380564 265294 380568
rect 265358 380566 265406 380626
rect 270953 380624 271006 380628
rect 271070 380626 271076 380628
rect 270953 380568 270958 380624
rect 265358 380564 265364 380566
rect 270953 380564 271006 380568
rect 271070 380566 271110 380626
rect 408677 380624 408702 380628
rect 408766 380626 408772 380628
rect 413456 380626 413462 380628
rect 408677 380568 408682 380624
rect 271070 380564 271076 380566
rect 408677 380564 408702 380568
rect 408766 380566 408834 380626
rect 413370 380566 413462 380626
rect 408766 380564 408772 380566
rect 413456 380564 413462 380566
rect 413526 380564 413532 380628
rect 419440 380564 419446 380628
rect 419510 380626 419516 380628
rect 419510 380566 419598 380626
rect 434345 380624 434406 380628
rect 434345 380568 434350 380624
rect 419510 380564 419516 380566
rect 434345 380564 434406 380568
rect 434470 380626 434476 380628
rect 434470 380566 434502 380626
rect 445937 380624 445966 380628
rect 446030 380626 446036 380628
rect 445937 380568 445942 380624
rect 434470 380564 434476 380566
rect 445937 380564 445966 380568
rect 446030 380566 446094 380626
rect 446030 380564 446036 380566
rect 254485 380563 254551 380564
rect 255865 380563 255931 380564
rect 256969 380563 257035 380564
rect 259453 380563 259519 380564
rect 260672 380490 260732 380564
rect 265249 380563 265315 380564
rect 270953 380563 271019 380564
rect 408677 380563 408743 380564
rect 413461 380563 413527 380564
rect 419441 380563 419507 380564
rect 434345 380563 434411 380564
rect 445937 380563 446003 380564
rect 253890 380430 260732 380490
rect 217060 380428 217066 380430
rect 203057 380354 203123 380357
rect 212809 380354 212875 380357
rect 213729 380354 213795 380357
rect 200070 380352 213795 380354
rect 200070 380296 203062 380352
rect 203118 380296 212814 380352
rect 212870 380296 213734 380352
rect 213790 380296 213795 380352
rect 200070 380294 213795 380296
rect 128353 380291 128419 380292
rect 155953 380291 156019 380292
rect 203057 380291 203123 380294
rect 212809 380291 212875 380294
rect 213729 380291 213795 380294
rect 119102 380156 119108 380220
rect 119172 380218 119178 380220
rect 208117 380218 208183 380221
rect 119172 380216 208183 380218
rect 119172 380160 208122 380216
rect 208178 380160 208183 380216
rect 119172 380158 208183 380160
rect 119172 380156 119178 380158
rect 208117 380155 208183 380158
rect 47577 380082 47643 380085
rect 217133 380082 217199 380085
rect 47577 380080 217199 380082
rect 47577 380024 47582 380080
rect 47638 380024 217138 380080
rect 217194 380024 217199 380080
rect 47577 380022 217199 380024
rect 47577 380019 47643 380022
rect 217133 380019 217199 380022
rect 216673 379674 216739 379677
rect 217869 379674 217935 379677
rect 216673 379672 217935 379674
rect 216673 379616 216678 379672
rect 216734 379616 217874 379672
rect 217930 379616 217935 379672
rect 216673 379614 217935 379616
rect 216673 379611 216739 379614
rect 217869 379611 217935 379614
rect 50286 379476 50292 379540
rect 50356 379538 50362 379540
rect 50981 379538 51047 379541
rect 50356 379536 51047 379538
rect 50356 379480 50986 379536
rect 51042 379480 51047 379536
rect 50356 379478 51047 379480
rect 50356 379476 50362 379478
rect 50981 379475 51047 379478
rect 202638 379476 202644 379540
rect 202708 379538 202714 379540
rect 202781 379538 202847 379541
rect 202708 379536 202847 379538
rect 202708 379480 202786 379536
rect 202842 379480 202847 379536
rect 202708 379478 202847 379480
rect 202708 379476 202714 379478
rect 202781 379475 202847 379478
rect 209078 379476 209084 379540
rect 209148 379538 209154 379540
rect 209589 379538 209655 379541
rect 209148 379536 209655 379538
rect 209148 379480 209594 379536
rect 209650 379480 209655 379536
rect 209148 379478 209655 379480
rect 209148 379476 209154 379478
rect 209589 379475 209655 379478
rect 217133 379538 217199 379541
rect 217685 379538 217751 379541
rect 217133 379536 217751 379538
rect 217133 379480 217138 379536
rect 217194 379480 217690 379536
rect 217746 379480 217751 379536
rect 217133 379478 217751 379480
rect 217133 379475 217199 379478
rect 217685 379475 217751 379478
rect 364374 379476 364380 379540
rect 364444 379538 364450 379540
rect 365621 379538 365687 379541
rect 364444 379536 365687 379538
rect 364444 379480 365626 379536
rect 365682 379480 365687 379536
rect 364444 379478 365687 379480
rect 364444 379476 364450 379478
rect 365621 379475 365687 379478
rect 47761 379402 47827 379405
rect 85481 379404 85547 379405
rect 86585 379404 86651 379405
rect 87689 379404 87755 379405
rect 79542 379402 79548 379404
rect 47761 379400 79548 379402
rect 47761 379344 47766 379400
rect 47822 379344 79548 379400
rect 47761 379342 79548 379344
rect 47761 379339 47827 379342
rect 79542 379340 79548 379342
rect 79612 379340 79618 379404
rect 85430 379402 85436 379404
rect 85390 379342 85436 379402
rect 85500 379400 85547 379404
rect 86534 379402 86540 379404
rect 85542 379344 85547 379400
rect 85430 379340 85436 379342
rect 85500 379340 85547 379344
rect 86494 379342 86540 379402
rect 86604 379400 86651 379404
rect 87638 379402 87644 379404
rect 86646 379344 86651 379400
rect 86534 379340 86540 379342
rect 86604 379340 86651 379344
rect 87598 379342 87644 379402
rect 87708 379400 87755 379404
rect 87750 379344 87755 379400
rect 87638 379340 87644 379342
rect 87708 379340 87755 379344
rect 85481 379339 85547 379340
rect 86585 379339 86651 379340
rect 87689 379339 87755 379340
rect 88333 379404 88399 379405
rect 88793 379404 88859 379405
rect 90081 379404 90147 379405
rect 88333 379400 88380 379404
rect 88444 379402 88450 379404
rect 88742 379402 88748 379404
rect 88333 379344 88338 379400
rect 88333 379340 88380 379344
rect 88444 379342 88490 379402
rect 88702 379342 88748 379402
rect 88812 379400 88859 379404
rect 90030 379402 90036 379404
rect 88854 379344 88859 379400
rect 88444 379340 88450 379342
rect 88742 379340 88748 379342
rect 88812 379340 88859 379344
rect 89990 379342 90036 379402
rect 90100 379400 90147 379404
rect 90142 379344 90147 379400
rect 90030 379340 90036 379342
rect 90100 379340 90147 379344
rect 88333 379339 88399 379340
rect 88793 379339 88859 379340
rect 90081 379339 90147 379340
rect 90633 379402 90699 379405
rect 91369 379404 91435 379405
rect 90766 379402 90772 379404
rect 90633 379400 90772 379402
rect 90633 379344 90638 379400
rect 90694 379344 90772 379400
rect 90633 379342 90772 379344
rect 90633 379339 90699 379342
rect 90766 379340 90772 379342
rect 90836 379340 90842 379404
rect 91318 379402 91324 379404
rect 91278 379342 91324 379402
rect 91388 379400 91435 379404
rect 91430 379344 91435 379400
rect 91318 379340 91324 379342
rect 91388 379340 91435 379344
rect 91369 379339 91435 379340
rect 92381 379404 92447 379405
rect 93485 379404 93551 379405
rect 96061 379404 96127 379405
rect 92381 379400 92428 379404
rect 92492 379402 92498 379404
rect 92381 379344 92386 379400
rect 92381 379340 92428 379344
rect 92492 379342 92538 379402
rect 93485 379400 93532 379404
rect 93596 379402 93602 379404
rect 93485 379344 93490 379400
rect 92492 379340 92498 379342
rect 93485 379340 93532 379344
rect 93596 379342 93642 379402
rect 96061 379400 96108 379404
rect 96172 379402 96178 379404
rect 96061 379344 96066 379400
rect 93596 379340 93602 379342
rect 96061 379340 96108 379344
rect 96172 379342 96218 379402
rect 96172 379340 96178 379342
rect 98126 379340 98132 379404
rect 98196 379402 98202 379404
rect 98269 379402 98335 379405
rect 98196 379400 98335 379402
rect 98196 379344 98274 379400
rect 98330 379344 98335 379400
rect 98196 379342 98335 379344
rect 98196 379340 98202 379342
rect 92381 379339 92447 379340
rect 93485 379339 93551 379340
rect 96061 379339 96127 379340
rect 98269 379339 98335 379342
rect 98453 379404 98519 379405
rect 101029 379404 101095 379405
rect 98453 379400 98500 379404
rect 98564 379402 98570 379404
rect 98453 379344 98458 379400
rect 98453 379340 98500 379344
rect 98564 379342 98610 379402
rect 101029 379400 101076 379404
rect 101140 379402 101146 379404
rect 101029 379344 101034 379400
rect 98564 379340 98570 379342
rect 101029 379340 101076 379344
rect 101140 379342 101186 379402
rect 101140 379340 101146 379342
rect 103278 379340 103284 379404
rect 103348 379402 103354 379404
rect 103513 379402 103579 379405
rect 103348 379400 103579 379402
rect 103348 379344 103518 379400
rect 103574 379344 103579 379400
rect 103348 379342 103579 379344
rect 103348 379340 103354 379342
rect 98453 379339 98519 379340
rect 101029 379339 101095 379340
rect 103513 379339 103579 379342
rect 105261 379402 105327 379405
rect 108205 379404 108271 379405
rect 108849 379404 108915 379405
rect 111241 379404 111307 379405
rect 105854 379402 105860 379404
rect 105261 379400 105860 379402
rect 105261 379344 105266 379400
rect 105322 379344 105860 379400
rect 105261 379342 105860 379344
rect 105261 379339 105327 379342
rect 105854 379340 105860 379342
rect 105924 379340 105930 379404
rect 108205 379400 108252 379404
rect 108316 379402 108322 379404
rect 108798 379402 108804 379404
rect 108205 379344 108210 379400
rect 108205 379340 108252 379344
rect 108316 379342 108362 379402
rect 108758 379342 108804 379402
rect 108868 379400 108915 379404
rect 111190 379402 111196 379404
rect 108910 379344 108915 379400
rect 108316 379340 108322 379342
rect 108798 379340 108804 379342
rect 108868 379340 108915 379344
rect 111150 379342 111196 379402
rect 111260 379400 111307 379404
rect 111302 379344 111307 379400
rect 111190 379340 111196 379342
rect 111260 379340 111307 379344
rect 112294 379340 112300 379404
rect 112364 379402 112370 379404
rect 112621 379402 112687 379405
rect 113449 379404 113515 379405
rect 113398 379402 113404 379404
rect 112364 379400 112687 379402
rect 112364 379344 112626 379400
rect 112682 379344 112687 379400
rect 112364 379342 112687 379344
rect 113358 379342 113404 379402
rect 113468 379400 113515 379404
rect 113510 379344 113515 379400
rect 112364 379340 112370 379342
rect 108205 379339 108271 379340
rect 108849 379339 108915 379340
rect 111241 379339 111307 379340
rect 112621 379339 112687 379342
rect 113398 379340 113404 379342
rect 113468 379340 113515 379344
rect 113449 379339 113515 379340
rect 114461 379404 114527 379405
rect 117129 379404 117195 379405
rect 141049 379404 141115 379405
rect 148593 379404 148659 379405
rect 150985 379404 151051 379405
rect 153561 379404 153627 379405
rect 183185 379404 183251 379405
rect 114461 379400 114508 379404
rect 114572 379402 114578 379404
rect 117078 379402 117084 379404
rect 114461 379344 114466 379400
rect 114461 379340 114508 379344
rect 114572 379342 114618 379402
rect 117038 379342 117084 379402
rect 117148 379400 117195 379404
rect 140998 379402 141004 379404
rect 117190 379344 117195 379400
rect 114572 379340 114578 379342
rect 117078 379340 117084 379342
rect 117148 379340 117195 379344
rect 140958 379342 141004 379402
rect 141068 379400 141115 379404
rect 148542 379402 148548 379404
rect 141110 379344 141115 379400
rect 140998 379340 141004 379342
rect 141068 379340 141115 379344
rect 148502 379342 148548 379402
rect 148612 379400 148659 379404
rect 150934 379402 150940 379404
rect 148654 379344 148659 379400
rect 148542 379340 148548 379342
rect 148612 379340 148659 379344
rect 150894 379342 150940 379402
rect 151004 379400 151051 379404
rect 153510 379402 153516 379404
rect 151046 379344 151051 379400
rect 150934 379340 150940 379342
rect 151004 379340 151051 379344
rect 153470 379342 153516 379402
rect 153580 379400 153627 379404
rect 183134 379402 183140 379404
rect 153622 379344 153627 379400
rect 153510 379340 153516 379342
rect 153580 379340 153627 379344
rect 183094 379342 183140 379402
rect 183204 379400 183251 379404
rect 183246 379344 183251 379400
rect 183134 379340 183140 379342
rect 183204 379340 183251 379344
rect 114461 379339 114527 379340
rect 117129 379339 117195 379340
rect 141049 379339 141115 379340
rect 148593 379339 148659 379340
rect 150985 379339 151051 379340
rect 153561 379339 153627 379340
rect 183185 379339 183251 379340
rect 199009 379402 199075 379405
rect 199510 379402 199516 379404
rect 199009 379400 199516 379402
rect 199009 379344 199014 379400
rect 199070 379344 199516 379400
rect 199009 379342 199516 379344
rect 199009 379339 199075 379342
rect 199510 379340 199516 379342
rect 199580 379340 199586 379404
rect 246021 379402 246087 379405
rect 247493 379404 247559 379405
rect 248597 379404 248663 379405
rect 250069 379404 250135 379405
rect 251173 379404 251239 379405
rect 252277 379404 252343 379405
rect 253381 379404 253447 379405
rect 246430 379402 246436 379404
rect 246021 379400 246436 379402
rect 246021 379344 246026 379400
rect 246082 379344 246436 379400
rect 246021 379342 246436 379344
rect 246021 379339 246087 379342
rect 246430 379340 246436 379342
rect 246500 379340 246506 379404
rect 247493 379400 247540 379404
rect 247604 379402 247610 379404
rect 247493 379344 247498 379400
rect 247493 379340 247540 379344
rect 247604 379342 247650 379402
rect 248597 379400 248644 379404
rect 248708 379402 248714 379404
rect 248597 379344 248602 379400
rect 247604 379340 247610 379342
rect 248597 379340 248644 379344
rect 248708 379342 248754 379402
rect 250069 379400 250116 379404
rect 250180 379402 250186 379404
rect 250069 379344 250074 379400
rect 248708 379340 248714 379342
rect 250069 379340 250116 379344
rect 250180 379342 250226 379402
rect 251173 379400 251220 379404
rect 251284 379402 251290 379404
rect 251173 379344 251178 379400
rect 250180 379340 250186 379342
rect 251173 379340 251220 379344
rect 251284 379342 251330 379402
rect 252277 379400 252324 379404
rect 252388 379402 252394 379404
rect 252277 379344 252282 379400
rect 251284 379340 251290 379342
rect 252277 379340 252324 379344
rect 252388 379342 252434 379402
rect 253381 379400 253428 379404
rect 253492 379402 253498 379404
rect 253381 379344 253386 379400
rect 252388 379340 252394 379342
rect 253381 379340 253428 379344
rect 253492 379342 253538 379402
rect 253492 379340 253498 379342
rect 257838 379340 257844 379404
rect 257908 379402 257914 379404
rect 258073 379402 258139 379405
rect 257908 379400 258139 379402
rect 257908 379344 258078 379400
rect 258134 379344 258139 379400
rect 257908 379342 258139 379344
rect 257908 379340 257914 379342
rect 247493 379339 247559 379340
rect 248597 379339 248663 379340
rect 250069 379339 250135 379340
rect 251173 379339 251239 379340
rect 252277 379339 252343 379340
rect 253381 379339 253447 379340
rect 258073 379339 258139 379342
rect 261661 379404 261727 379405
rect 268653 379404 268719 379405
rect 271045 379404 271111 379405
rect 261661 379400 261708 379404
rect 261772 379402 261778 379404
rect 261661 379344 261666 379400
rect 261661 379340 261708 379344
rect 261772 379342 261818 379402
rect 268653 379400 268700 379404
rect 268764 379402 268770 379404
rect 268653 379344 268658 379400
rect 261772 379340 261778 379342
rect 268653 379340 268700 379344
rect 268764 379342 268810 379402
rect 271045 379400 271092 379404
rect 271156 379402 271162 379404
rect 272057 379402 272123 379405
rect 273253 379404 273319 379405
rect 272190 379402 272196 379404
rect 271045 379344 271050 379400
rect 268764 379340 268770 379342
rect 271045 379340 271092 379344
rect 271156 379342 271202 379402
rect 272057 379400 272196 379402
rect 272057 379344 272062 379400
rect 272118 379344 272196 379400
rect 272057 379342 272196 379344
rect 271156 379340 271162 379342
rect 261661 379339 261727 379340
rect 268653 379339 268719 379340
rect 271045 379339 271111 379340
rect 272057 379339 272123 379342
rect 272190 379340 272196 379342
rect 272260 379340 272266 379404
rect 273253 379400 273300 379404
rect 273364 379402 273370 379404
rect 274173 379402 274239 379405
rect 275645 379404 275711 379405
rect 276013 379404 276079 379405
rect 276933 379404 276999 379405
rect 285949 379404 286015 379405
rect 274398 379402 274404 379404
rect 273253 379344 273258 379400
rect 273253 379340 273300 379344
rect 273364 379342 273410 379402
rect 274173 379400 274404 379402
rect 274173 379344 274178 379400
rect 274234 379344 274404 379400
rect 274173 379342 274404 379344
rect 273364 379340 273370 379342
rect 273253 379339 273319 379340
rect 274173 379339 274239 379342
rect 274398 379340 274404 379342
rect 274468 379340 274474 379404
rect 275645 379400 275692 379404
rect 275756 379402 275762 379404
rect 275645 379344 275650 379400
rect 275645 379340 275692 379344
rect 275756 379342 275802 379402
rect 276013 379400 276060 379404
rect 276124 379402 276130 379404
rect 276013 379344 276018 379400
rect 275756 379340 275762 379342
rect 276013 379340 276060 379344
rect 276124 379342 276170 379402
rect 276933 379400 276980 379404
rect 277044 379402 277050 379404
rect 278078 379402 278084 379404
rect 276933 379344 276938 379400
rect 276124 379340 276130 379342
rect 276933 379340 276980 379344
rect 277044 379342 277090 379402
rect 277902 379342 278084 379402
rect 277044 379340 277050 379342
rect 275645 379339 275711 379340
rect 276013 379339 276079 379340
rect 276933 379339 276999 379340
rect 277902 379269 277962 379342
rect 278078 379340 278084 379342
rect 278148 379340 278154 379404
rect 285949 379400 285996 379404
rect 286060 379402 286066 379404
rect 287697 379402 287763 379405
rect 290917 379404 290983 379405
rect 288198 379402 288204 379404
rect 285949 379344 285954 379400
rect 285949 379340 285996 379344
rect 286060 379342 286106 379402
rect 287697 379400 288204 379402
rect 287697 379344 287702 379400
rect 287758 379344 288204 379400
rect 287697 379342 288204 379344
rect 286060 379340 286066 379342
rect 285949 379339 286015 379340
rect 287697 379339 287763 379342
rect 288198 379340 288204 379342
rect 288268 379340 288274 379404
rect 290917 379400 290964 379404
rect 291028 379402 291034 379404
rect 292665 379402 292731 379405
rect 295885 379404 295951 379405
rect 298461 379404 298527 379405
rect 300853 379404 300919 379405
rect 293350 379402 293356 379404
rect 290917 379344 290922 379400
rect 290917 379340 290964 379344
rect 291028 379342 291074 379402
rect 292665 379400 293356 379402
rect 292665 379344 292670 379400
rect 292726 379344 293356 379400
rect 292665 379342 293356 379344
rect 291028 379340 291034 379342
rect 290917 379339 290983 379340
rect 292665 379339 292731 379342
rect 293350 379340 293356 379342
rect 293420 379340 293426 379404
rect 295885 379400 295932 379404
rect 295996 379402 296002 379404
rect 295885 379344 295890 379400
rect 295885 379340 295932 379344
rect 295996 379342 296042 379402
rect 298461 379400 298508 379404
rect 298572 379402 298578 379404
rect 298461 379344 298466 379400
rect 295996 379340 296002 379342
rect 298461 379340 298508 379344
rect 298572 379342 298618 379402
rect 300853 379400 300900 379404
rect 300964 379402 300970 379404
rect 302785 379402 302851 379405
rect 305821 379404 305887 379405
rect 310973 379404 311039 379405
rect 313365 379404 313431 379405
rect 315757 379404 315823 379405
rect 303470 379402 303476 379404
rect 300853 379344 300858 379400
rect 298572 379340 298578 379342
rect 300853 379340 300900 379344
rect 300964 379342 301010 379402
rect 302785 379400 303476 379402
rect 302785 379344 302790 379400
rect 302846 379344 303476 379400
rect 302785 379342 303476 379344
rect 300964 379340 300970 379342
rect 295885 379339 295951 379340
rect 298461 379339 298527 379340
rect 300853 379339 300919 379340
rect 302785 379339 302851 379342
rect 303470 379340 303476 379342
rect 303540 379340 303546 379404
rect 305821 379400 305868 379404
rect 305932 379402 305938 379404
rect 305821 379344 305826 379400
rect 305821 379340 305868 379344
rect 305932 379342 305978 379402
rect 310973 379400 311020 379404
rect 311084 379402 311090 379404
rect 310973 379344 310978 379400
rect 305932 379340 305938 379342
rect 310973 379340 311020 379344
rect 311084 379342 311130 379402
rect 313365 379400 313412 379404
rect 313476 379402 313482 379404
rect 313365 379344 313370 379400
rect 311084 379340 311090 379342
rect 313365 379340 313412 379344
rect 313476 379342 313522 379402
rect 315757 379400 315804 379404
rect 315868 379402 315874 379404
rect 317413 379402 317479 379405
rect 323301 379404 323367 379405
rect 325969 379404 326035 379405
rect 343449 379404 343515 379405
rect 396073 379404 396139 379405
rect 318374 379402 318380 379404
rect 315757 379344 315762 379400
rect 313476 379340 313482 379342
rect 315757 379340 315804 379344
rect 315868 379342 315914 379402
rect 317413 379400 318380 379402
rect 317413 379344 317418 379400
rect 317474 379344 318380 379400
rect 317413 379342 318380 379344
rect 315868 379340 315874 379342
rect 305821 379339 305887 379340
rect 310973 379339 311039 379340
rect 313365 379339 313431 379340
rect 315757 379339 315823 379340
rect 317413 379339 317479 379342
rect 318374 379340 318380 379342
rect 318444 379340 318450 379404
rect 323301 379400 323348 379404
rect 323412 379402 323418 379404
rect 325918 379402 325924 379404
rect 323301 379344 323306 379400
rect 323301 379340 323348 379344
rect 323412 379342 323458 379402
rect 325878 379342 325924 379402
rect 325988 379400 326035 379404
rect 343398 379402 343404 379404
rect 326030 379344 326035 379400
rect 323412 379340 323418 379342
rect 325918 379340 325924 379342
rect 325988 379340 326035 379344
rect 343358 379342 343404 379402
rect 343468 379400 343515 379404
rect 396022 379402 396028 379404
rect 343510 379344 343515 379400
rect 343398 379340 343404 379342
rect 343468 379340 343515 379344
rect 395982 379342 396028 379402
rect 396092 379400 396139 379404
rect 396134 379344 396139 379400
rect 396022 379340 396028 379342
rect 396092 379340 396139 379344
rect 323301 379339 323367 379340
rect 325969 379339 326035 379340
rect 343449 379339 343515 379340
rect 396073 379339 396139 379340
rect 397085 379404 397151 379405
rect 397085 379400 397132 379404
rect 397196 379402 397202 379404
rect 403617 379402 403683 379405
rect 404118 379402 404124 379404
rect 397085 379344 397090 379400
rect 397085 379340 397132 379344
rect 397196 379342 397242 379402
rect 403617 379400 404124 379402
rect 403617 379344 403622 379400
rect 403678 379344 404124 379400
rect 403617 379342 404124 379344
rect 397196 379340 397202 379342
rect 397085 379339 397151 379340
rect 403617 379339 403683 379342
rect 404118 379340 404124 379342
rect 404188 379340 404194 379404
rect 405825 379402 405891 379405
rect 407573 379404 407639 379405
rect 408309 379404 408375 379405
rect 411253 379404 411319 379405
rect 412357 379404 412423 379405
rect 406510 379402 406516 379404
rect 405825 379400 406516 379402
rect 405825 379344 405830 379400
rect 405886 379344 406516 379400
rect 405825 379342 406516 379344
rect 405825 379339 405891 379342
rect 406510 379340 406516 379342
rect 406580 379340 406586 379404
rect 407573 379400 407620 379404
rect 407684 379402 407690 379404
rect 407573 379344 407578 379400
rect 407573 379340 407620 379344
rect 407684 379342 407730 379402
rect 408309 379400 408356 379404
rect 408420 379402 408426 379404
rect 408309 379344 408314 379400
rect 407684 379340 407690 379342
rect 408309 379340 408356 379344
rect 408420 379342 408466 379402
rect 411253 379400 411300 379404
rect 411364 379402 411370 379404
rect 411253 379344 411258 379400
rect 408420 379340 408426 379342
rect 411253 379340 411300 379344
rect 411364 379342 411410 379402
rect 412357 379400 412404 379404
rect 412468 379402 412474 379404
rect 413093 379402 413159 379405
rect 414565 379404 414631 379405
rect 423397 379404 423463 379405
rect 426433 379404 426499 379405
rect 413502 379402 413508 379404
rect 412357 379344 412362 379400
rect 411364 379340 411370 379342
rect 412357 379340 412404 379344
rect 412468 379342 412514 379402
rect 413093 379400 413508 379402
rect 413093 379344 413098 379400
rect 413154 379344 413508 379400
rect 413093 379342 413508 379344
rect 412468 379340 412474 379342
rect 407573 379339 407639 379340
rect 408309 379339 408375 379340
rect 411253 379339 411319 379340
rect 412357 379339 412423 379340
rect 413093 379339 413159 379342
rect 413502 379340 413508 379342
rect 413572 379340 413578 379404
rect 414565 379400 414612 379404
rect 414676 379402 414682 379404
rect 414565 379344 414570 379400
rect 414565 379340 414612 379344
rect 414676 379342 414722 379402
rect 423397 379400 423444 379404
rect 423508 379402 423514 379404
rect 426382 379402 426388 379404
rect 423397 379344 423402 379400
rect 414676 379340 414682 379342
rect 423397 379340 423444 379344
rect 423508 379342 423554 379402
rect 426342 379342 426388 379402
rect 426452 379400 426499 379404
rect 426494 379344 426499 379400
rect 423508 379340 423514 379342
rect 426382 379340 426388 379342
rect 426452 379340 426499 379344
rect 414565 379339 414631 379340
rect 423397 379339 423463 379340
rect 426433 379339 426499 379340
rect 426617 379402 426683 379405
rect 435725 379404 435791 379405
rect 439037 379404 439103 379405
rect 427486 379402 427492 379404
rect 426617 379400 427492 379402
rect 426617 379344 426622 379400
rect 426678 379344 427492 379400
rect 426617 379342 427492 379344
rect 426617 379339 426683 379342
rect 427486 379340 427492 379342
rect 427556 379340 427562 379404
rect 435725 379400 435772 379404
rect 435836 379402 435842 379404
rect 435725 379344 435730 379400
rect 435725 379340 435772 379344
rect 435836 379342 435882 379402
rect 439037 379400 439084 379404
rect 439148 379402 439154 379404
rect 447501 379402 447567 379405
rect 450997 379404 451063 379405
rect 448278 379402 448284 379404
rect 439037 379344 439042 379400
rect 435836 379340 435842 379342
rect 439037 379340 439084 379344
rect 439148 379342 439194 379402
rect 447501 379400 448284 379402
rect 447501 379344 447506 379400
rect 447562 379344 448284 379400
rect 447501 379342 448284 379344
rect 439148 379340 439154 379342
rect 435725 379339 435791 379340
rect 439037 379339 439103 379340
rect 447501 379339 447567 379342
rect 448278 379340 448284 379342
rect 448348 379340 448354 379404
rect 450997 379400 451044 379404
rect 451108 379402 451114 379404
rect 452745 379402 452811 379405
rect 453430 379402 453436 379404
rect 450997 379344 451002 379400
rect 450997 379340 451044 379344
rect 451108 379342 451154 379402
rect 452745 379400 453436 379402
rect 452745 379344 452750 379400
rect 452806 379344 453436 379400
rect 452745 379342 453436 379344
rect 451108 379340 451114 379342
rect 450997 379339 451063 379340
rect 452745 379339 452811 379342
rect 453430 379340 453436 379342
rect 453500 379340 453506 379404
rect 455597 379402 455663 379405
rect 458357 379404 458423 379405
rect 460933 379404 460999 379405
rect 463509 379404 463575 379405
rect 455822 379402 455828 379404
rect 455597 379400 455828 379402
rect 455597 379344 455602 379400
rect 455658 379344 455828 379400
rect 455597 379342 455828 379344
rect 455597 379339 455663 379342
rect 455822 379340 455828 379342
rect 455892 379340 455898 379404
rect 458357 379400 458404 379404
rect 458468 379402 458474 379404
rect 458357 379344 458362 379400
rect 458357 379340 458404 379344
rect 458468 379342 458514 379402
rect 460933 379400 460980 379404
rect 461044 379402 461050 379404
rect 460933 379344 460938 379400
rect 458468 379340 458474 379342
rect 460933 379340 460980 379344
rect 461044 379342 461090 379402
rect 463509 379400 463556 379404
rect 463620 379402 463626 379404
rect 474825 379402 474891 379405
rect 475878 379402 475884 379404
rect 463509 379344 463514 379400
rect 461044 379340 461050 379342
rect 463509 379340 463556 379344
rect 463620 379342 463666 379402
rect 474825 379400 475884 379402
rect 474825 379344 474830 379400
rect 474886 379344 475884 379400
rect 474825 379342 475884 379344
rect 463620 379340 463626 379342
rect 458357 379339 458423 379340
rect 460933 379339 460999 379340
rect 463509 379339 463575 379340
rect 474825 379339 474891 379342
rect 475878 379340 475884 379342
rect 475948 379340 475954 379404
rect 47669 379266 47735 379269
rect 80421 379268 80487 379269
rect 78254 379266 78260 379268
rect 47669 379264 78260 379266
rect 47669 379208 47674 379264
rect 47730 379208 78260 379264
rect 47669 379206 78260 379208
rect 47669 379203 47735 379206
rect 78254 379204 78260 379206
rect 78324 379204 78330 379268
rect 80421 379264 80468 379268
rect 80532 379266 80538 379268
rect 81433 379266 81499 379269
rect 95969 379268 96035 379269
rect 99465 379268 99531 379269
rect 102961 379268 103027 379269
rect 81750 379266 81756 379268
rect 80421 379208 80426 379264
rect 80421 379204 80468 379208
rect 80532 379206 80578 379266
rect 81433 379264 81756 379266
rect 81433 379208 81438 379264
rect 81494 379208 81756 379264
rect 81433 379206 81756 379208
rect 80532 379204 80538 379206
rect 80421 379203 80487 379204
rect 81433 379203 81499 379206
rect 81750 379204 81756 379206
rect 81820 379266 81826 379268
rect 95918 379266 95924 379268
rect 81820 379206 93870 379266
rect 95878 379206 95924 379266
rect 95988 379264 96035 379268
rect 99414 379266 99420 379268
rect 96030 379208 96035 379264
rect 81820 379204 81826 379206
rect 79542 379068 79548 379132
rect 79612 379130 79618 379132
rect 93810 379130 93870 379206
rect 95918 379204 95924 379206
rect 95988 379204 96035 379208
rect 99374 379206 99420 379266
rect 99484 379264 99531 379268
rect 102910 379266 102916 379268
rect 99526 379208 99531 379264
rect 99414 379204 99420 379206
rect 99484 379204 99531 379208
rect 102870 379206 102916 379266
rect 102980 379264 103027 379268
rect 103022 379208 103027 379264
rect 102910 379204 102916 379206
rect 102980 379204 103027 379208
rect 105302 379204 105308 379268
rect 105372 379266 105378 379268
rect 105537 379266 105603 379269
rect 105372 379264 105603 379266
rect 105372 379208 105542 379264
rect 105598 379208 105603 379264
rect 105372 379206 105603 379208
rect 105372 379204 105378 379206
rect 95969 379203 96035 379204
rect 99465 379203 99531 379204
rect 102961 379203 103027 379204
rect 105537 379203 105603 379206
rect 109718 379204 109724 379268
rect 109788 379266 109794 379268
rect 213821 379266 213887 379269
rect 277853 379266 277962 379269
rect 109788 379206 211354 379266
rect 109788 379204 109794 379206
rect 207565 379130 207631 379133
rect 207933 379130 207999 379133
rect 79612 379070 85682 379130
rect 93810 379128 207999 379130
rect 93810 379072 207570 379128
rect 207626 379072 207938 379128
rect 207994 379072 207999 379128
rect 93810 379070 207999 379072
rect 211294 379130 211354 379206
rect 213821 379264 277962 379266
rect 213821 379208 213826 379264
rect 213882 379208 277858 379264
rect 277914 379208 277962 379264
rect 213821 379206 277962 379208
rect 278037 379266 278103 379269
rect 279141 379268 279207 379269
rect 278446 379266 278452 379268
rect 278037 379264 278452 379266
rect 278037 379208 278042 379264
rect 278098 379208 278452 379264
rect 278037 379206 278452 379208
rect 213821 379203 213887 379206
rect 277853 379203 277919 379206
rect 278037 379203 278103 379206
rect 278446 379204 278452 379206
rect 278516 379204 278522 379268
rect 279141 379264 279188 379268
rect 279252 379266 279258 379268
rect 280705 379266 280771 379269
rect 280838 379266 280844 379268
rect 279141 379208 279146 379264
rect 279141 379204 279188 379208
rect 279252 379206 279298 379266
rect 280705 379264 280844 379266
rect 280705 379208 280710 379264
rect 280766 379208 280844 379264
rect 280705 379206 280844 379208
rect 279252 379204 279258 379206
rect 279141 379203 279207 379204
rect 280705 379203 280771 379206
rect 280838 379204 280844 379206
rect 280908 379204 280914 379268
rect 283005 379266 283071 379269
rect 283414 379266 283420 379268
rect 283005 379264 283420 379266
rect 283005 379208 283010 379264
rect 283066 379208 283420 379264
rect 283005 379206 283420 379208
rect 283005 379203 283071 379206
rect 283414 379204 283420 379206
rect 283484 379204 283490 379268
rect 371141 379266 371207 379269
rect 402973 379268 403039 379269
rect 405365 379268 405431 379269
rect 398230 379266 398236 379268
rect 371141 379264 398236 379266
rect 371141 379208 371146 379264
rect 371202 379208 398236 379264
rect 371141 379206 398236 379208
rect 371141 379203 371207 379206
rect 398230 379204 398236 379206
rect 398300 379204 398306 379268
rect 402973 379264 403020 379268
rect 403084 379266 403090 379268
rect 402973 379208 402978 379264
rect 402973 379204 403020 379208
rect 403084 379206 403130 379266
rect 405365 379264 405412 379268
rect 405476 379266 405482 379268
rect 410057 379266 410123 379269
rect 410742 379266 410748 379268
rect 405365 379208 405370 379264
rect 403084 379204 403090 379206
rect 405365 379204 405412 379208
rect 405476 379206 405522 379266
rect 410057 379264 410748 379266
rect 410057 379208 410062 379264
rect 410118 379208 410748 379264
rect 410057 379206 410748 379208
rect 405476 379204 405482 379206
rect 402973 379203 403039 379204
rect 405365 379203 405431 379204
rect 410057 379203 410123 379206
rect 410742 379204 410748 379206
rect 410812 379204 410818 379268
rect 415761 379266 415827 379269
rect 416037 379268 416103 379269
rect 415894 379266 415900 379268
rect 415761 379264 415900 379266
rect 415761 379208 415766 379264
rect 415822 379208 415900 379264
rect 415761 379206 415900 379208
rect 415761 379203 415827 379206
rect 415894 379204 415900 379206
rect 415964 379204 415970 379268
rect 416037 379264 416084 379268
rect 416148 379266 416154 379268
rect 437749 379266 437815 379269
rect 473445 379268 473511 379269
rect 437974 379266 437980 379268
rect 416037 379208 416042 379264
rect 416037 379204 416084 379208
rect 416148 379206 416194 379266
rect 437749 379264 437980 379266
rect 437749 379208 437754 379264
rect 437810 379208 437980 379264
rect 437749 379206 437980 379208
rect 416148 379204 416154 379206
rect 416037 379203 416103 379204
rect 437749 379203 437815 379206
rect 437974 379204 437980 379206
rect 438044 379204 438050 379268
rect 473445 379264 473492 379268
rect 473556 379266 473562 379268
rect 480529 379266 480595 379269
rect 503069 379268 503135 379269
rect 503529 379268 503595 379269
rect 480846 379266 480852 379268
rect 473445 379208 473450 379264
rect 473445 379204 473492 379208
rect 473556 379206 473602 379266
rect 480529 379264 480852 379266
rect 480529 379208 480534 379264
rect 480590 379208 480852 379264
rect 480529 379206 480852 379208
rect 473556 379204 473562 379206
rect 473445 379203 473511 379204
rect 480529 379203 480595 379206
rect 480846 379204 480852 379206
rect 480916 379204 480922 379268
rect 503069 379264 503116 379268
rect 503180 379266 503186 379268
rect 503069 379208 503074 379264
rect 503069 379204 503116 379208
rect 503180 379206 503226 379266
rect 503180 379204 503186 379206
rect 503478 379204 503484 379268
rect 503548 379266 503595 379268
rect 503548 379264 503640 379266
rect 503590 379208 503640 379264
rect 503548 379206 503640 379208
rect 503548 379204 503595 379206
rect 503069 379203 503135 379204
rect 503529 379203 503595 379204
rect 211705 379130 211771 379133
rect 218329 379130 218395 379133
rect 239254 379130 239260 379132
rect 211294 379128 218395 379130
rect 211294 379072 211710 379128
rect 211766 379072 218334 379128
rect 218390 379072 218395 379128
rect 211294 379070 218395 379072
rect 79612 379068 79618 379070
rect 47577 378994 47643 378997
rect 47761 378994 47827 378997
rect 47577 378992 47827 378994
rect 47577 378936 47582 378992
rect 47638 378936 47766 378992
rect 47822 378936 47827 378992
rect 47577 378934 47827 378936
rect 47577 378931 47643 378934
rect 47761 378931 47827 378934
rect 78254 378932 78260 378996
rect 78324 378994 78330 378996
rect 85622 378994 85682 379070
rect 207565 379067 207631 379070
rect 207933 379067 207999 379070
rect 211705 379067 211771 379070
rect 218329 379067 218395 379070
rect 238710 379070 239260 379130
rect 208853 378994 208919 378997
rect 238710 378994 238770 379070
rect 239254 379068 239260 379070
rect 239324 379130 239330 379132
rect 365529 379130 365595 379133
rect 399518 379130 399524 379132
rect 239324 379128 399524 379130
rect 239324 379072 365534 379128
rect 365590 379072 399524 379128
rect 239324 379070 399524 379072
rect 239324 379068 239330 379070
rect 365529 379067 365595 379070
rect 399518 379068 399524 379070
rect 399588 379068 399594 379132
rect 433374 379130 433380 379132
rect 412590 379070 433380 379130
rect 78324 378934 84210 378994
rect 85622 378992 238770 378994
rect 85622 378936 208858 378992
rect 208914 378936 238770 378992
rect 85622 378934 238770 378936
rect 78324 378932 78330 378934
rect 43989 378860 44055 378861
rect 43989 378858 44036 378860
rect 43944 378856 44036 378858
rect 43944 378800 43994 378856
rect 43944 378798 44036 378800
rect 43989 378796 44036 378798
rect 44100 378796 44106 378860
rect 83222 378796 83228 378860
rect 83292 378858 83298 378860
rect 83457 378858 83523 378861
rect 83292 378856 83523 378858
rect 83292 378800 83462 378856
rect 83518 378800 83523 378856
rect 83292 378798 83523 378800
rect 84150 378858 84210 378934
rect 208853 378931 208919 378934
rect 241462 378932 241468 378996
rect 241532 378994 241538 378996
rect 373165 378994 373231 378997
rect 241532 378992 373231 378994
rect 241532 378936 373170 378992
rect 373226 378936 373231 378992
rect 241532 378934 373231 378936
rect 241532 378932 241538 378934
rect 373165 378931 373231 378934
rect 376886 378932 376892 378996
rect 376956 378994 376962 378996
rect 412590 378994 412650 379070
rect 433374 379068 433380 379070
rect 433444 379068 433450 379132
rect 465073 379130 465139 379133
rect 465942 379130 465948 379132
rect 465073 379128 465948 379130
rect 465073 379072 465078 379128
rect 465134 379072 465948 379128
rect 465073 379070 465948 379072
rect 465073 379067 465139 379070
rect 465942 379068 465948 379070
rect 466012 379068 466018 379132
rect 376956 378934 412650 378994
rect 477585 378994 477651 378997
rect 483381 378996 483447 378997
rect 478454 378994 478460 378996
rect 477585 378992 478460 378994
rect 477585 378936 477590 378992
rect 477646 378936 478460 378992
rect 477585 378934 478460 378936
rect 376956 378932 376962 378934
rect 477585 378931 477651 378934
rect 478454 378932 478460 378934
rect 478524 378932 478530 378996
rect 483381 378992 483428 378996
rect 483492 378994 483498 378996
rect 483381 378936 483386 378992
rect 483381 378932 483428 378936
rect 483492 378934 483538 378994
rect 483492 378932 483498 378934
rect 483381 378931 483447 378932
rect 207933 378858 207999 378861
rect 248229 378860 248295 378861
rect 241830 378858 241836 378860
rect 84150 378798 200130 378858
rect 83292 378796 83298 378798
rect 43989 378795 44055 378796
rect 83457 378795 83523 378798
rect 94681 378724 94747 378725
rect 94630 378722 94636 378724
rect 94590 378662 94636 378722
rect 94700 378720 94747 378724
rect 94742 378664 94747 378720
rect 94630 378660 94636 378662
rect 94700 378660 94747 378664
rect 97022 378660 97028 378724
rect 97092 378722 97098 378724
rect 97165 378722 97231 378725
rect 138473 378724 138539 378725
rect 138422 378722 138428 378724
rect 97092 378720 97231 378722
rect 97092 378664 97170 378720
rect 97226 378664 97231 378720
rect 97092 378662 97231 378664
rect 138382 378662 138428 378722
rect 138492 378720 138539 378724
rect 138534 378664 138539 378720
rect 97092 378660 97098 378662
rect 94681 378659 94747 378660
rect 97165 378659 97231 378662
rect 138422 378660 138428 378662
rect 138492 378660 138539 378664
rect 200070 378722 200130 378798
rect 207933 378856 241836 378858
rect 207933 378800 207938 378856
rect 207994 378800 241836 378856
rect 207933 378798 241836 378800
rect 207933 378795 207999 378798
rect 241830 378796 241836 378798
rect 241900 378796 241906 378860
rect 248229 378856 248276 378860
rect 248340 378858 248346 378860
rect 252369 378858 252435 378861
rect 375005 378858 375071 378861
rect 402278 378858 402284 378860
rect 248229 378800 248234 378856
rect 248229 378796 248276 378800
rect 248340 378798 248386 378858
rect 252369 378856 402284 378858
rect 252369 378800 252374 378856
rect 252430 378800 375010 378856
rect 375066 378800 402284 378856
rect 252369 378798 402284 378800
rect 248340 378796 248346 378798
rect 248229 378795 248295 378796
rect 252369 378795 252435 378798
rect 375005 378795 375071 378798
rect 402278 378796 402284 378798
rect 402348 378796 402354 378860
rect 467925 378858 467991 378861
rect 470869 378860 470935 378861
rect 468518 378858 468524 378860
rect 467925 378856 468524 378858
rect 467925 378800 467930 378856
rect 467986 378800 468524 378856
rect 467925 378798 468524 378800
rect 467925 378795 467991 378798
rect 468518 378796 468524 378798
rect 468588 378796 468594 378860
rect 470869 378856 470916 378860
rect 470980 378858 470986 378860
rect 470869 378800 470874 378856
rect 470869 378796 470916 378800
rect 470980 378798 471026 378858
rect 470980 378796 470986 378798
rect 470869 378795 470935 378796
rect 208209 378722 208275 378725
rect 238150 378722 238156 378724
rect 200070 378720 238156 378722
rect 200070 378664 208214 378720
rect 208270 378664 238156 378720
rect 200070 378662 238156 378664
rect 138473 378659 138539 378660
rect 208209 378659 208275 378662
rect 238150 378660 238156 378662
rect 238220 378722 238226 378724
rect 371141 378722 371207 378725
rect 238220 378720 371207 378722
rect 238220 378664 371146 378720
rect 371202 378664 371207 378720
rect 238220 378662 371207 378664
rect 238220 378660 238226 378662
rect 371141 378659 371207 378662
rect 373165 378722 373231 378725
rect 400438 378722 400444 378724
rect 373165 378720 400444 378722
rect 373165 378664 373170 378720
rect 373226 378664 400444 378720
rect 373165 378662 400444 378664
rect 373165 378659 373231 378662
rect 400438 378660 400444 378662
rect 400508 378660 400514 378724
rect 418245 378722 418311 378725
rect 425973 378724 426039 378725
rect 418470 378722 418476 378724
rect 418245 378720 418476 378722
rect 418245 378664 418250 378720
rect 418306 378664 418476 378720
rect 418245 378662 418476 378664
rect 418245 378659 418311 378662
rect 418470 378660 418476 378662
rect 418540 378660 418546 378724
rect 425973 378720 426020 378724
rect 426084 378722 426090 378724
rect 427905 378722 427971 378725
rect 428222 378722 428228 378724
rect 425973 378664 425978 378720
rect 425973 378660 426020 378664
rect 426084 378662 426130 378722
rect 427905 378720 428228 378722
rect 427905 378664 427910 378720
rect 427966 378664 428228 378720
rect 427905 378662 428228 378664
rect 426084 378660 426090 378662
rect 425973 378659 426039 378660
rect 427905 378659 427971 378662
rect 428222 378660 428228 378662
rect 428292 378660 428298 378724
rect 115790 378524 115796 378588
rect 115860 378586 115866 378588
rect 206829 378586 206895 378589
rect 212625 378586 212691 378589
rect 115860 378584 212691 378586
rect 115860 378528 206834 378584
rect 206890 378528 212630 378584
rect 212686 378528 212691 378584
rect 115860 378526 212691 378528
rect 115860 378524 115866 378526
rect 206829 378523 206895 378526
rect 212625 378523 212691 378526
rect 218329 378586 218395 378589
rect 253565 378588 253631 378589
rect 258349 378588 258415 378589
rect 260925 378588 260991 378589
rect 263593 378588 263659 378589
rect 218329 378584 253306 378586
rect 218329 378528 218334 378584
rect 218390 378528 253306 378584
rect 218329 378526 253306 378528
rect 218329 378523 218395 378526
rect 80421 378450 80487 378453
rect 221089 378450 221155 378453
rect 240542 378450 240548 378452
rect 80421 378448 240548 378450
rect 80421 378392 80426 378448
rect 80482 378392 221094 378448
rect 221150 378392 240548 378448
rect 80421 378390 240548 378392
rect 80421 378387 80487 378390
rect 221089 378387 221155 378390
rect 240542 378388 240548 378390
rect 240612 378450 240618 378452
rect 241462 378450 241468 378452
rect 240612 378390 241468 378450
rect 240612 378388 240618 378390
rect 241462 378388 241468 378390
rect 241532 378388 241538 378452
rect 241830 378388 241836 378452
rect 241900 378450 241906 378452
rect 252369 378450 252435 378453
rect 241900 378448 252435 378450
rect 241900 378392 252374 378448
rect 252430 378392 252435 378448
rect 241900 378390 252435 378392
rect 253246 378450 253306 378526
rect 253565 378584 253612 378588
rect 253676 378586 253682 378588
rect 253565 378528 253570 378584
rect 253565 378524 253612 378528
rect 253676 378526 253722 378586
rect 258349 378584 258396 378588
rect 258460 378586 258466 378588
rect 258349 378528 258354 378584
rect 253676 378524 253682 378526
rect 258349 378524 258396 378528
rect 258460 378526 258506 378586
rect 260925 378584 260972 378588
rect 261036 378586 261042 378588
rect 263542 378586 263548 378588
rect 260925 378528 260930 378584
rect 258460 378524 258466 378526
rect 260925 378524 260972 378528
rect 261036 378526 261082 378586
rect 263502 378526 263548 378586
rect 263612 378584 263659 378588
rect 263654 378528 263659 378584
rect 261036 378524 261042 378526
rect 263542 378524 263548 378526
rect 263612 378524 263659 378528
rect 253565 378523 253631 378524
rect 258349 378523 258415 378524
rect 260925 378523 260991 378524
rect 263593 378523 263659 378524
rect 265893 378588 265959 378589
rect 265893 378584 265940 378588
rect 266004 378586 266010 378588
rect 268101 378586 268167 378589
rect 273437 378588 273503 378589
rect 320909 378588 320975 378589
rect 416957 378588 417023 378589
rect 268326 378586 268332 378588
rect 265893 378528 265898 378584
rect 265893 378524 265940 378528
rect 266004 378526 266050 378586
rect 268101 378584 268332 378586
rect 268101 378528 268106 378584
rect 268162 378528 268332 378584
rect 268101 378526 268332 378528
rect 266004 378524 266010 378526
rect 265893 378523 265959 378524
rect 268101 378523 268167 378526
rect 268326 378524 268332 378526
rect 268396 378524 268402 378588
rect 273437 378584 273484 378588
rect 273548 378586 273554 378588
rect 273437 378528 273442 378584
rect 273437 378524 273484 378528
rect 273548 378526 273594 378586
rect 320909 378584 320956 378588
rect 321020 378586 321026 378588
rect 320909 378528 320914 378584
rect 273548 378524 273554 378526
rect 320909 378524 320956 378528
rect 321020 378526 321066 378586
rect 416957 378584 417004 378588
rect 417068 378586 417074 378588
rect 436461 378586 436527 378589
rect 436870 378586 436876 378588
rect 416957 378528 416962 378584
rect 321020 378524 321026 378526
rect 416957 378524 417004 378528
rect 417068 378526 417114 378586
rect 436461 378584 436876 378586
rect 436461 378528 436466 378584
rect 436522 378528 436876 378584
rect 436461 378526 436876 378528
rect 417068 378524 417074 378526
rect 273437 378523 273503 378524
rect 320909 378523 320975 378524
rect 416957 378523 417023 378524
rect 436461 378523 436527 378526
rect 436870 378524 436876 378526
rect 436940 378524 436946 378588
rect 262857 378450 262923 378453
rect 253246 378448 262923 378450
rect 253246 378392 262862 378448
rect 262918 378392 262923 378448
rect 253246 378390 262923 378392
rect 241900 378388 241906 378390
rect 252369 378387 252435 378390
rect 262857 378387 262923 378390
rect 343173 378452 343239 378453
rect 343173 378448 343220 378452
rect 343284 378450 343290 378452
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 343173 378392 343178 378448
rect 343173 378388 343220 378392
rect 343284 378390 343330 378450
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 343284 378388 343290 378390
rect 343173 378387 343239 378388
rect 580165 378387 580231 378390
rect 104014 378252 104020 378316
rect 104084 378314 104090 378316
rect 104433 378314 104499 378317
rect 107561 378316 107627 378317
rect 107510 378314 107516 378316
rect 104084 378312 104499 378314
rect 104084 378256 104438 378312
rect 104494 378256 104499 378312
rect 104084 378254 104499 378256
rect 107470 378254 107516 378314
rect 107580 378312 107627 378316
rect 107622 378256 107627 378312
rect 104084 378252 104090 378254
rect 104433 378251 104499 378254
rect 107510 378252 107516 378254
rect 107580 378252 107627 378256
rect 118182 378252 118188 378316
rect 118252 378314 118258 378316
rect 213821 378314 213887 378317
rect 244273 378316 244339 378317
rect 244222 378314 244228 378316
rect 118252 378312 213887 378314
rect 118252 378256 213826 378312
rect 213882 378256 213887 378312
rect 118252 378254 213887 378256
rect 244182 378254 244228 378314
rect 244292 378312 244339 378316
rect 244334 378256 244339 378312
rect 118252 378252 118258 378254
rect 107561 378251 107627 378252
rect 213821 378251 213887 378254
rect 244222 378252 244228 378254
rect 244292 378252 244339 378256
rect 244273 378251 244339 378252
rect 250621 378316 250687 378317
rect 262765 378316 262831 378317
rect 266353 378316 266419 378317
rect 250621 378312 250668 378316
rect 250732 378314 250738 378316
rect 250621 378256 250626 378312
rect 250621 378252 250668 378256
rect 250732 378254 250778 378314
rect 262765 378312 262812 378316
rect 262876 378314 262882 378316
rect 266302 378314 266308 378316
rect 262765 378256 262770 378312
rect 250732 378252 250738 378254
rect 262765 378252 262812 378256
rect 262876 378254 262922 378314
rect 266262 378254 266308 378314
rect 266372 378312 266419 378316
rect 266414 378256 266419 378312
rect 262876 378252 262882 378254
rect 266302 378252 266308 378254
rect 266372 378252 266419 378256
rect 250621 378251 250687 378252
rect 262765 378251 262831 378252
rect 266353 378251 266419 378252
rect 267549 378316 267615 378317
rect 431125 378316 431191 378317
rect 267549 378312 267596 378316
rect 267660 378314 267666 378316
rect 267549 378256 267554 378312
rect 267549 378252 267596 378256
rect 267660 378254 267706 378314
rect 431125 378312 431172 378316
rect 431236 378314 431242 378316
rect 431125 378256 431130 378312
rect 267660 378252 267666 378254
rect 431125 378252 431172 378256
rect 431236 378254 431282 378314
rect 583520 378300 584960 378390
rect 431236 378252 431242 378254
rect 267549 378251 267615 378252
rect 431125 378251 431191 378252
rect 84326 378116 84332 378180
rect 84396 378178 84402 378180
rect 85021 378178 85087 378181
rect 101857 378180 101923 378181
rect 106457 378180 106523 378181
rect 84396 378176 85087 378178
rect 84396 378120 85026 378176
rect 85082 378120 85087 378176
rect 84396 378118 85087 378120
rect 84396 378116 84402 378118
rect 85021 378115 85087 378118
rect 100702 378116 100708 378180
rect 100772 378116 100778 378180
rect 101806 378178 101812 378180
rect 101766 378118 101812 378178
rect 101876 378176 101923 378180
rect 106406 378178 106412 378180
rect 101918 378120 101923 378176
rect 101806 378116 101812 378118
rect 101876 378116 101923 378120
rect 106366 378118 106412 378178
rect 106476 378176 106523 378180
rect 106518 378120 106523 378176
rect 106406 378116 106412 378118
rect 106476 378116 106523 378120
rect 100710 378042 100770 378116
rect 101857 378115 101923 378116
rect 106457 378115 106523 378116
rect 182265 378178 182331 378181
rect 182817 378178 182883 378181
rect 183502 378178 183508 378180
rect 182265 378176 183508 378178
rect 182265 378120 182270 378176
rect 182326 378120 182822 378176
rect 182878 378120 183508 378176
rect 182265 378118 183508 378120
rect 182265 378115 182331 378118
rect 182817 378115 182883 378118
rect 183502 378116 183508 378118
rect 183572 378116 183578 378180
rect 211654 378116 211660 378180
rect 211724 378178 211730 378180
rect 212441 378178 212507 378181
rect 211724 378176 212507 378178
rect 211724 378120 212446 378176
rect 212502 378120 212507 378176
rect 211724 378118 212507 378120
rect 211724 378116 211730 378118
rect 212441 378115 212507 378118
rect 212625 378178 212691 378181
rect 274633 378178 274699 378181
rect 212625 378176 274699 378178
rect 212625 378120 212630 378176
rect 212686 378120 274638 378176
rect 274694 378120 274699 378176
rect 212625 378118 274699 378120
rect 212625 378115 212691 378118
rect 274633 378115 274699 378118
rect 308622 378116 308628 378180
rect 308692 378116 308698 378180
rect 371601 378178 371667 378181
rect 409965 378180 410031 378181
rect 418153 378180 418219 378181
rect 376886 378178 376892 378180
rect 371601 378176 376892 378178
rect 371601 378120 371606 378176
rect 371662 378120 376892 378176
rect 371601 378118 376892 378120
rect 100710 377982 200130 378042
rect 199142 377844 199148 377908
rect 199212 377906 199218 377908
rect 199469 377906 199535 377909
rect 199212 377904 199535 377906
rect 199212 377848 199474 377904
rect 199530 377848 199535 377904
rect 199212 377846 199535 377848
rect 200070 377906 200130 377982
rect 217542 377980 217548 378044
rect 217612 378042 217618 378044
rect 308630 378042 308690 378116
rect 371601 378115 371667 378118
rect 376886 378116 376892 378118
rect 376956 378116 376962 378180
rect 409965 378176 410012 378180
rect 410076 378178 410082 378180
rect 418102 378178 418108 378180
rect 409965 378120 409970 378176
rect 409965 378116 410012 378120
rect 410076 378118 410122 378178
rect 418062 378118 418108 378178
rect 418172 378176 418219 378180
rect 418214 378120 418219 378176
rect 410076 378116 410082 378118
rect 418102 378116 418108 378118
rect 418172 378116 418219 378120
rect 409965 378115 410031 378116
rect 418153 378115 418219 378116
rect 419625 378178 419691 378181
rect 421741 378180 421807 378181
rect 423949 378180 424015 378181
rect 420678 378178 420684 378180
rect 419625 378176 420684 378178
rect 419625 378120 419630 378176
rect 419686 378120 420684 378176
rect 419625 378118 420684 378120
rect 419625 378115 419691 378118
rect 420678 378116 420684 378118
rect 420748 378116 420754 378180
rect 421741 378176 421788 378180
rect 421852 378178 421858 378180
rect 421741 378120 421746 378176
rect 421741 378116 421788 378120
rect 421852 378118 421898 378178
rect 423949 378176 423996 378180
rect 424060 378178 424066 378180
rect 425145 378178 425211 378181
rect 425278 378178 425284 378180
rect 423949 378120 423954 378176
rect 421852 378116 421858 378118
rect 423949 378116 423996 378120
rect 424060 378118 424106 378178
rect 425145 378176 425284 378178
rect 425145 378120 425150 378176
rect 425206 378120 425284 378176
rect 425145 378118 425284 378120
rect 424060 378116 424066 378118
rect 421741 378115 421807 378116
rect 423949 378115 424015 378116
rect 425145 378115 425211 378118
rect 425278 378116 425284 378118
rect 425348 378116 425354 378180
rect 428273 378178 428339 378181
rect 428590 378178 428596 378180
rect 428273 378176 428596 378178
rect 428273 378120 428278 378176
rect 428334 378120 428596 378176
rect 428273 378118 428596 378120
rect 428273 378115 428339 378118
rect 428590 378116 428596 378118
rect 428660 378116 428666 378180
rect 429285 378178 429351 378181
rect 432229 378180 432295 378181
rect 429694 378178 429700 378180
rect 429285 378176 429700 378178
rect 429285 378120 429290 378176
rect 429346 378120 429700 378176
rect 429285 378118 429700 378120
rect 429285 378115 429351 378118
rect 429694 378116 429700 378118
rect 429764 378116 429770 378180
rect 432229 378176 432276 378180
rect 432340 378178 432346 378180
rect 432229 378120 432234 378176
rect 432229 378116 432276 378120
rect 432340 378118 432386 378178
rect 432340 378116 432346 378118
rect 432229 378115 432295 378116
rect 217612 377982 308690 378042
rect 217612 377980 217618 377982
rect 359774 377980 359780 378044
rect 359844 378042 359850 378044
rect 463509 378042 463575 378045
rect 359844 378040 463575 378042
rect 359844 377984 463514 378040
rect 463570 377984 463575 378040
rect 359844 377982 463575 377984
rect 359844 377980 359850 377982
rect 463509 377979 463575 377982
rect 216622 377906 216628 377908
rect 200070 377846 216628 377906
rect 199212 377844 199218 377846
rect 199469 377843 199535 377846
rect 216622 377844 216628 377846
rect 216692 377906 216698 377908
rect 217409 377906 217475 377909
rect 216692 377904 217475 377906
rect 216692 377848 217414 377904
rect 217470 377848 217475 377904
rect 216692 377846 217475 377848
rect 216692 377844 216698 377846
rect 217409 377843 217475 377846
rect 213678 376756 213684 376820
rect 213748 376818 213754 376820
rect 213821 376818 213887 376821
rect 213748 376816 213887 376818
rect 213748 376760 213826 376816
rect 213882 376760 213887 376816
rect 213748 376758 213887 376760
rect 213748 376756 213754 376758
rect 213821 376755 213887 376758
rect 370078 376756 370084 376820
rect 370148 376818 370154 376820
rect 371141 376818 371207 376821
rect 370148 376816 371207 376818
rect 370148 376760 371146 376816
rect 371202 376760 371207 376816
rect 370148 376758 371207 376760
rect 370148 376756 370154 376758
rect 371141 376755 371207 376758
rect 377438 376620 377444 376684
rect 377508 376682 377514 376684
rect 483381 376682 483447 376685
rect 377508 376680 483447 376682
rect 377508 376624 483386 376680
rect 483442 376624 483447 376680
rect 377508 376622 483447 376624
rect 377508 376620 377514 376622
rect 483381 376619 483447 376622
rect 212625 376410 212691 376413
rect 213545 376410 213611 376413
rect 212625 376408 213611 376410
rect 212625 376352 212630 376408
rect 212686 376352 213550 376408
rect 213606 376352 213611 376408
rect 212625 376350 213611 376352
rect 212625 376347 212691 376350
rect 213545 376347 213611 376350
rect 209814 375532 209820 375596
rect 209884 375594 209890 375596
rect 210969 375594 211035 375597
rect 209884 375592 211035 375594
rect 209884 375536 210974 375592
rect 211030 375536 211035 375592
rect 209884 375534 211035 375536
rect 209884 375532 209890 375534
rect 210969 375531 211035 375534
rect 213862 375532 213868 375596
rect 213932 375594 213938 375596
rect 215109 375594 215175 375597
rect 213932 375592 215175 375594
rect 213932 375536 215114 375592
rect 215170 375536 215175 375592
rect 213932 375534 215175 375536
rect 213932 375532 213938 375534
rect 215109 375531 215175 375534
rect 54385 375458 54451 375461
rect 57094 375458 57100 375460
rect 54385 375456 57100 375458
rect 54385 375400 54390 375456
rect 54446 375400 57100 375456
rect 54385 375398 57100 375400
rect 54385 375395 54451 375398
rect 57094 375396 57100 375398
rect 57164 375396 57170 375460
rect 208894 375396 208900 375460
rect 208964 375458 208970 375460
rect 209497 375458 209563 375461
rect 208964 375456 209563 375458
rect 208964 375400 209502 375456
rect 209558 375400 209563 375456
rect 208964 375398 209563 375400
rect 208964 375396 208970 375398
rect 209497 375395 209563 375398
rect 209998 375396 210004 375460
rect 210068 375458 210074 375460
rect 211061 375458 211127 375461
rect 210068 375456 211127 375458
rect 210068 375400 211066 375456
rect 211122 375400 211127 375456
rect 210068 375398 211127 375400
rect 210068 375396 210074 375398
rect 211061 375395 211127 375398
rect 214046 375396 214052 375460
rect 214116 375458 214122 375460
rect 215201 375458 215267 375461
rect 214116 375456 215267 375458
rect 214116 375400 215206 375456
rect 215262 375400 215267 375456
rect 214116 375398 215267 375400
rect 214116 375396 214122 375398
rect 215201 375395 215267 375398
rect 377438 375260 377444 375324
rect 377508 375322 377514 375324
rect 379605 375322 379671 375325
rect 377508 375320 379671 375322
rect 377508 375264 379610 375320
rect 379666 375264 379671 375320
rect 377508 375262 379671 375264
rect 377508 375260 377514 375262
rect 379605 375259 379671 375262
rect 375414 375124 375420 375188
rect 375484 375186 375490 375188
rect 376661 375186 376727 375189
rect 375484 375184 376727 375186
rect 375484 375128 376666 375184
rect 376722 375128 376727 375184
rect 375484 375126 376727 375128
rect 375484 375124 375490 375126
rect 376661 375123 376727 375126
rect 217501 374916 217567 374917
rect 217501 374912 217548 374916
rect 217612 374914 217618 374916
rect 217501 374856 217506 374912
rect 217501 374852 217548 374856
rect 217612 374854 217658 374914
rect 217612 374852 217618 374854
rect 217501 374851 217567 374852
rect 377949 374780 378015 374781
rect 377949 374776 377996 374780
rect 378060 374778 378066 374780
rect 377949 374720 377954 374776
rect 377949 374716 377996 374720
rect 378060 374718 378106 374778
rect 378060 374716 378066 374718
rect 377949 374715 378015 374716
rect 199377 371924 199443 371925
rect 199326 371922 199332 371924
rect 199250 371862 199332 371922
rect 199396 371922 199443 371924
rect 359733 371922 359799 371925
rect 359917 371922 359983 371925
rect 199396 371920 359983 371922
rect 199438 371864 359738 371920
rect 359794 371864 359922 371920
rect 359978 371864 359983 371920
rect 199326 371860 199332 371862
rect 199396 371862 359983 371864
rect 199396 371860 199443 371862
rect 199377 371859 199443 371860
rect 359733 371859 359799 371862
rect 359917 371859 359983 371862
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect 178534 358804 178540 358868
rect 178604 358866 178610 358868
rect 178677 358866 178743 358869
rect 178604 358864 178743 358866
rect 178604 358808 178682 358864
rect 178738 358808 178743 358864
rect 178604 358806 178743 358808
rect 178604 358804 178610 358806
rect 178677 358803 178743 358806
rect 179638 358804 179644 358868
rect 179708 358866 179714 358868
rect 179873 358866 179939 358869
rect 190913 358868 190979 358869
rect 338481 358868 338547 358869
rect 190862 358866 190868 358868
rect 179708 358864 179939 358866
rect 179708 358808 179878 358864
rect 179934 358808 179939 358864
rect 179708 358806 179939 358808
rect 190822 358806 190868 358866
rect 190932 358864 190979 358868
rect 338430 358866 338436 358868
rect 190974 358808 190979 358864
rect 179708 358804 179714 358806
rect 179873 358803 179939 358806
rect 190862 358804 190868 358806
rect 190932 358804 190979 358808
rect 338390 358806 338436 358866
rect 338500 358864 338547 358868
rect 338542 358808 338547 358864
rect 338430 358804 338436 358806
rect 338500 358804 338547 358808
rect 339718 358804 339724 358868
rect 339788 358866 339794 358868
rect 339861 358866 339927 358869
rect 339788 358864 339927 358866
rect 339788 358808 339866 358864
rect 339922 358808 339927 358864
rect 339788 358806 339927 358808
rect 339788 358804 339794 358806
rect 190913 358803 190979 358804
rect 338481 358803 338547 358804
rect 339861 358803 339927 358806
rect 350942 358804 350948 358868
rect 351012 358866 351018 358868
rect 351729 358866 351795 358869
rect 351012 358864 351795 358866
rect 351012 358808 351734 358864
rect 351790 358808 351795 358864
rect 351012 358806 351795 358808
rect 351012 358804 351018 358806
rect 351729 358803 351795 358806
rect 498510 358804 498516 358868
rect 498580 358866 498586 358868
rect 498929 358866 498995 358869
rect 498580 358864 498995 358866
rect 498580 358808 498934 358864
rect 498990 358808 498995 358864
rect 498580 358806 498995 358808
rect 498580 358804 498586 358806
rect 498929 358803 498995 358806
rect 499798 358804 499804 358868
rect 499868 358866 499874 358868
rect 500769 358866 500835 358869
rect 510889 358868 510955 358869
rect 510838 358866 510844 358868
rect 499868 358864 500835 358866
rect 499868 358808 500774 358864
rect 500830 358808 500835 358864
rect 499868 358806 500835 358808
rect 510798 358806 510844 358866
rect 510908 358864 510955 358868
rect 510950 358808 510955 358864
rect 499868 358804 499874 358806
rect 500769 358803 500835 358806
rect 510838 358804 510844 358806
rect 510908 358804 510955 358808
rect 510889 358803 510955 358804
rect -960 358458 480 358548
rect 3601 358458 3667 358461
rect -960 358456 3667 358458
rect -960 358400 3606 358456
rect 3662 358400 3667 358456
rect -960 358398 3667 358400
rect -960 358308 480 358398
rect 3601 358395 3667 358398
rect 196558 353154 196618 353190
rect 198825 353154 198891 353157
rect 196558 353152 198891 353154
rect 196558 353096 198830 353152
rect 198886 353096 198891 353152
rect 196558 353094 198891 353096
rect 356562 353154 356622 353190
rect 358905 353154 358971 353157
rect 356562 353152 358971 353154
rect 356562 353096 358910 353152
rect 358966 353096 358971 353152
rect 356562 353094 358971 353096
rect 198825 353091 198891 353094
rect 358905 353091 358971 353094
rect 516558 353018 516618 353190
rect 519077 353018 519143 353021
rect 519445 353018 519511 353021
rect 516558 353016 519511 353018
rect 516558 352960 519082 353016
rect 519138 352960 519450 353016
rect 519506 352960 519511 353016
rect 516558 352958 519511 352960
rect 519077 352955 519143 352958
rect 519445 352955 519511 352958
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect 57513 311130 57579 311133
rect 57513 311128 60062 311130
rect 57513 311072 57518 311128
rect 57574 311072 60062 311128
rect 57513 311070 60062 311072
rect 57513 311067 57579 311070
rect 60002 310894 60062 311070
rect 217501 310994 217567 310997
rect 376937 310994 377003 310997
rect 217501 310992 219450 310994
rect 217501 310936 217506 310992
rect 217562 310936 219450 310992
rect 217501 310934 219450 310936
rect 217501 310931 217567 310934
rect 219390 310924 219450 310934
rect 376937 310992 379898 310994
rect 376937 310936 376942 310992
rect 376998 310936 379898 310992
rect 376937 310934 379898 310936
rect 376937 310931 377003 310934
rect 379838 310924 379898 310934
rect 219390 310864 220064 310924
rect 379838 310864 380052 310924
rect 57329 310450 57395 310453
rect 57789 310450 57855 310453
rect 57329 310448 60062 310450
rect 57329 310392 57334 310448
rect 57390 310392 57794 310448
rect 57850 310392 60062 310448
rect 57329 310390 60062 310392
rect 57329 310387 57395 310390
rect 57789 310387 57855 310390
rect 60002 309942 60062 310390
rect 217133 310042 217199 310045
rect 217961 310042 218027 310045
rect 377305 310042 377371 310045
rect 377857 310042 377923 310045
rect 217133 310040 219450 310042
rect 217133 309984 217138 310040
rect 217194 309984 217966 310040
rect 218022 309984 219450 310040
rect 217133 309982 219450 309984
rect 217133 309979 217199 309982
rect 217961 309979 218027 309982
rect 219390 309972 219450 309982
rect 377305 310040 379898 310042
rect 377305 309984 377310 310040
rect 377366 309984 377862 310040
rect 377918 309984 379898 310040
rect 377305 309982 379898 309984
rect 377305 309979 377371 309982
rect 377857 309979 377923 309982
rect 379838 309972 379898 309982
rect 219390 309912 220064 309972
rect 379838 309912 380052 309972
rect 56869 309090 56935 309093
rect 57697 309090 57763 309093
rect 56869 309088 57763 309090
rect 56869 309032 56874 309088
rect 56930 309032 57702 309088
rect 57758 309032 57763 309088
rect 56869 309030 57763 309032
rect 56869 309027 56935 309030
rect 57697 309027 57763 309030
rect 56869 307866 56935 307869
rect 217685 307866 217751 307869
rect 377673 307866 377739 307869
rect 56869 307864 59922 307866
rect 56869 307808 56874 307864
rect 56930 307808 59922 307864
rect 56869 307806 59922 307808
rect 56869 307803 56935 307806
rect 59862 307796 59922 307806
rect 217685 307864 219450 307866
rect 217685 307808 217690 307864
rect 217746 307808 219450 307864
rect 217685 307806 219450 307808
rect 217685 307803 217751 307806
rect 219390 307796 219450 307806
rect 377673 307864 379898 307866
rect 377673 307808 377678 307864
rect 377734 307808 379898 307864
rect 377673 307806 379898 307808
rect 377673 307803 377739 307806
rect 379838 307796 379898 307806
rect 59862 307736 60032 307796
rect 219390 307736 220064 307796
rect 379838 307736 380052 307796
rect 56777 307730 56843 307733
rect 57789 307730 57855 307733
rect 56777 307728 57855 307730
rect 56777 307672 56782 307728
rect 56838 307672 57794 307728
rect 57850 307672 57855 307728
rect 56777 307670 57855 307672
rect 56777 307667 56843 307670
rect 57789 307667 57855 307670
rect 217041 307730 217107 307733
rect 217501 307730 217567 307733
rect 217041 307728 217567 307730
rect 217041 307672 217046 307728
rect 217102 307672 217506 307728
rect 217562 307672 217567 307728
rect 217041 307670 217567 307672
rect 217041 307667 217107 307670
rect 217501 307667 217567 307670
rect 57789 306778 57855 306781
rect 60002 306778 60062 306814
rect 219390 306784 220064 306844
rect 379838 306784 380052 306844
rect 57789 306776 60062 306778
rect 57789 306720 57794 306776
rect 57850 306720 60062 306776
rect 57789 306718 60062 306720
rect 217501 306778 217567 306781
rect 219390 306778 219450 306784
rect 217501 306776 219450 306778
rect 217501 306720 217506 306776
rect 217562 306720 219450 306776
rect 217501 306718 219450 306720
rect 377765 306778 377831 306781
rect 379838 306778 379898 306784
rect 377765 306776 379898 306778
rect 377765 306720 377770 306776
rect 377826 306720 379898 306776
rect 377765 306718 379898 306720
rect 57789 306715 57855 306718
rect 217501 306715 217567 306718
rect 377765 306715 377831 306718
rect -960 306234 480 306324
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 57697 305010 57763 305013
rect 60002 305010 60062 305046
rect 219390 305016 220064 305076
rect 379470 305016 380052 305076
rect 57697 305008 60062 305010
rect 57697 304952 57702 305008
rect 57758 304952 60062 305008
rect 57697 304950 60062 304952
rect 216765 305010 216831 305013
rect 217317 305010 217383 305013
rect 219390 305010 219450 305016
rect 216765 305008 219450 305010
rect 216765 304952 216770 305008
rect 216826 304952 217322 305008
rect 217378 304952 219450 305008
rect 216765 304950 219450 304952
rect 377581 305010 377647 305013
rect 377765 305010 377831 305013
rect 379470 305010 379530 305016
rect 377581 305008 379530 305010
rect 377581 304952 377586 305008
rect 377642 304952 377770 305008
rect 377826 304952 379530 305008
rect 377581 304950 379530 304952
rect 57697 304947 57763 304950
rect 216765 304947 216831 304950
rect 217317 304947 217383 304950
rect 377581 304947 377647 304950
rect 377765 304947 377831 304950
rect 57605 303650 57671 303653
rect 60002 303650 60062 303958
rect 219390 303928 220064 303988
rect 379838 303928 380052 303988
rect 217777 303922 217843 303925
rect 219390 303922 219450 303928
rect 217777 303920 219450 303922
rect 217777 303864 217782 303920
rect 217838 303864 219450 303920
rect 217777 303862 219450 303864
rect 377489 303922 377555 303925
rect 379838 303922 379898 303928
rect 377489 303920 379898 303922
rect 377489 303864 377494 303920
rect 377550 303864 379898 303920
rect 377489 303862 379898 303864
rect 217777 303859 217843 303862
rect 377489 303859 377555 303862
rect 57605 303648 60062 303650
rect 57605 303592 57610 303648
rect 57666 303592 60062 303648
rect 57605 303590 60062 303592
rect 57605 303587 57671 303590
rect 57421 301610 57487 301613
rect 60002 301610 60062 302190
rect 219390 302160 220064 302220
rect 379838 302160 380052 302220
rect 216949 302154 217015 302157
rect 219390 302154 219450 302160
rect 216949 302152 219450 302154
rect 216949 302096 216954 302152
rect 217010 302096 219450 302152
rect 216949 302094 219450 302096
rect 377121 302154 377187 302157
rect 378041 302154 378107 302157
rect 379838 302154 379898 302160
rect 377121 302152 379898 302154
rect 377121 302096 377126 302152
rect 377182 302096 378046 302152
rect 378102 302096 379898 302152
rect 377121 302094 379898 302096
rect 216949 302091 217015 302094
rect 377121 302091 377187 302094
rect 378041 302091 378107 302094
rect 57421 301608 60062 301610
rect 57421 301552 57426 301608
rect 57482 301552 60062 301608
rect 57421 301550 60062 301552
rect 57421 301547 57487 301550
rect 583520 298604 584960 298844
rect 519353 293858 519419 293861
rect 516558 293856 519419 293858
rect 516558 293800 519358 293856
rect 519414 293800 519419 293856
rect 516558 293798 519419 293800
rect 516558 293350 516618 293798
rect 519353 293795 519419 293798
rect -960 293028 480 293268
rect 196558 292770 196618 293350
rect 199193 292770 199259 292773
rect 199653 292770 199719 292773
rect 196558 292768 199719 292770
rect 196558 292712 199198 292768
rect 199254 292712 199658 292768
rect 199714 292712 199719 292768
rect 196558 292710 199719 292712
rect 356562 292770 356622 293350
rect 359273 292770 359339 292773
rect 359549 292770 359615 292773
rect 356562 292768 359615 292770
rect 356562 292712 359278 292768
rect 359334 292712 359554 292768
rect 359610 292712 359615 292768
rect 356562 292710 359615 292712
rect 199193 292707 199259 292710
rect 199653 292707 199719 292710
rect 359273 292707 359339 292710
rect 359549 292707 359615 292710
rect 518893 292498 518959 292501
rect 519445 292498 519511 292501
rect 516558 292496 519511 292498
rect 516558 292440 518898 292496
rect 518954 292440 519450 292496
rect 519506 292440 519511 292496
rect 516558 292438 519511 292440
rect 358813 291818 358879 291821
rect 359457 291818 359523 291821
rect 356562 291816 359523 291818
rect 356562 291760 358818 291816
rect 358874 291760 359462 291816
rect 359518 291760 359523 291816
rect 356562 291758 359523 291760
rect 356562 291718 356622 291758
rect 358813 291755 358879 291758
rect 359457 291755 359523 291758
rect 516558 291718 516618 292438
rect 518893 292435 518959 292438
rect 519445 292435 519511 292438
rect 196558 291682 196618 291718
rect 198917 291682 198983 291685
rect 199469 291682 199535 291685
rect 196558 291680 199535 291682
rect 196558 291624 198922 291680
rect 198978 291624 199474 291680
rect 199530 291624 199535 291680
rect 196558 291622 199535 291624
rect 198917 291619 198983 291622
rect 199469 291619 199535 291622
rect 198733 291002 198799 291005
rect 199745 291002 199811 291005
rect 359181 291002 359247 291005
rect 196558 291000 199811 291002
rect 196558 290944 198738 291000
rect 198794 290944 199750 291000
rect 199806 290944 199811 291000
rect 196558 290942 199811 290944
rect 196558 290358 196618 290942
rect 198733 290939 198799 290942
rect 199745 290939 199811 290942
rect 356562 291000 359247 291002
rect 356562 290944 359186 291000
rect 359242 290944 359247 291000
rect 356562 290942 359247 290944
rect 356562 290358 356622 290942
rect 359181 290939 359247 290942
rect 516558 290322 516618 290358
rect 518985 290322 519051 290325
rect 519537 290322 519603 290325
rect 516558 290320 519603 290322
rect 516558 290264 518990 290320
rect 519046 290264 519542 290320
rect 519598 290264 519603 290320
rect 516558 290262 519603 290264
rect 518985 290259 519051 290262
rect 519537 290259 519603 290262
rect 196558 288826 196618 288862
rect 199009 288826 199075 288829
rect 196558 288824 199075 288826
rect 196558 288768 199014 288824
rect 199070 288768 199075 288824
rect 196558 288766 199075 288768
rect 356562 288826 356622 288862
rect 359733 288826 359799 288829
rect 356562 288824 359799 288826
rect 356562 288768 359738 288824
rect 359794 288768 359799 288824
rect 356562 288766 359799 288768
rect 199009 288763 199075 288766
rect 359733 288763 359799 288766
rect 516558 288554 516618 288862
rect 519169 288554 519235 288557
rect 519629 288554 519695 288557
rect 520181 288554 520247 288557
rect 516558 288552 520247 288554
rect 516558 288496 519174 288552
rect 519230 288496 519634 288552
rect 519690 288496 520186 288552
rect 520242 288496 520247 288552
rect 516558 288494 520247 288496
rect 519169 288491 519235 288494
rect 519629 288491 519695 288494
rect 520181 288491 520247 288494
rect 199101 288418 199167 288421
rect 199561 288418 199627 288421
rect 199101 288416 199627 288418
rect 199101 288360 199106 288416
rect 199162 288360 199566 288416
rect 199622 288360 199627 288416
rect 199101 288358 199627 288360
rect 199101 288355 199167 288358
rect 199561 288355 199627 288358
rect 196558 287602 196618 287638
rect 199101 287602 199167 287605
rect 196558 287600 199167 287602
rect 196558 287544 199106 287600
rect 199162 287544 199167 287600
rect 196558 287542 199167 287544
rect 356562 287602 356622 287638
rect 359089 287602 359155 287605
rect 356562 287600 359155 287602
rect 356562 287544 359094 287600
rect 359150 287544 359155 287600
rect 356562 287542 359155 287544
rect 516558 287602 516618 287638
rect 519261 287602 519327 287605
rect 516558 287600 519327 287602
rect 516558 287544 519266 287600
rect 519322 287544 519327 287600
rect 516558 287542 519327 287544
rect 199101 287539 199167 287542
rect 359089 287539 359155 287542
rect 519261 287539 519327 287542
rect 583520 285276 584960 285516
rect 58709 284202 58775 284205
rect 58709 284200 60062 284202
rect 58709 284144 58714 284200
rect 58770 284144 60062 284200
rect 58709 284142 60062 284144
rect 58709 284139 58775 284142
rect 60002 283966 60062 284142
rect 216673 284066 216739 284069
rect 376937 284066 377003 284069
rect 216673 284064 219450 284066
rect 216673 284008 216678 284064
rect 216734 284008 219450 284064
rect 216673 284006 219450 284008
rect 216673 284003 216739 284006
rect 219390 283996 219450 284006
rect 376937 284064 379530 284066
rect 376937 284008 376942 284064
rect 376998 284008 379530 284064
rect 376937 284006 379530 284008
rect 376937 284003 377003 284006
rect 379470 283996 379530 284006
rect 219390 283936 220064 283996
rect 379470 283936 380052 283996
rect 57237 282570 57303 282573
rect 57881 282570 57947 282573
rect 57237 282568 60062 282570
rect 57237 282512 57242 282568
rect 57298 282512 57886 282568
rect 57942 282512 60062 282568
rect 57237 282510 60062 282512
rect 57237 282507 57303 282510
rect 57881 282507 57947 282510
rect 60002 282334 60062 282510
rect 219390 282304 220064 282364
rect 379470 282304 380052 282364
rect 54201 282298 54267 282301
rect 54702 282298 54708 282300
rect 54201 282296 54708 282298
rect 54201 282240 54206 282296
rect 54262 282240 54708 282296
rect 54201 282238 54708 282240
rect 54201 282235 54267 282238
rect 54702 282236 54708 282238
rect 54772 282236 54778 282300
rect 216673 282298 216739 282301
rect 219390 282298 219450 282304
rect 216673 282296 219450 282298
rect 216673 282240 216678 282296
rect 216734 282240 219450 282296
rect 216673 282238 219450 282240
rect 376937 282298 377003 282301
rect 379470 282298 379530 282304
rect 376937 282296 379530 282298
rect 376937 282240 376942 282296
rect 376998 282240 379530 282296
rect 376937 282238 379530 282240
rect 216673 282235 216739 282238
rect 376937 282235 377003 282238
rect 216857 282162 216923 282165
rect 376753 282162 376819 282165
rect 216857 282160 219450 282162
rect 216857 282104 216862 282160
rect 216918 282104 219450 282160
rect 216857 282102 219450 282104
rect 216857 282099 216923 282102
rect 219390 282092 219450 282102
rect 376753 282160 379530 282162
rect 376753 282104 376758 282160
rect 376814 282104 379530 282160
rect 376753 282102 379530 282104
rect 376753 282099 376819 282102
rect 379470 282092 379530 282102
rect 58801 282026 58867 282029
rect 60002 282026 60062 282062
rect 219390 282032 220064 282092
rect 379470 282032 380052 282092
rect 58801 282024 60062 282026
rect 58801 281968 58806 282024
rect 58862 281968 60062 282024
rect 58801 281966 60062 281968
rect 58801 281963 58867 281966
rect -960 279972 480 280212
rect 95969 273868 96035 273869
rect 113357 273868 113423 273869
rect 95904 273804 95910 273868
rect 95974 273866 96035 273868
rect 95974 273864 96066 273866
rect 96030 273808 96066 273864
rect 95974 273806 96066 273808
rect 95974 273804 96035 273806
rect 113312 273804 113318 273868
rect 113382 273866 113423 273868
rect 273161 273866 273227 273869
rect 274400 273866 274406 273868
rect 113382 273864 113474 273866
rect 113418 273808 113474 273864
rect 113382 273806 113474 273808
rect 273161 273864 274406 273866
rect 273161 273808 273166 273864
rect 273222 273808 274406 273864
rect 273161 273806 274406 273808
rect 113382 273804 113423 273806
rect 95969 273803 96035 273804
rect 113357 273803 113423 273804
rect 273161 273803 273227 273806
rect 274400 273804 274406 273806
rect 274470 273804 274476 273868
rect 133413 273732 133479 273733
rect 133413 273730 133446 273732
rect 133354 273728 133446 273730
rect 133354 273672 133418 273728
rect 133354 273670 133446 273672
rect 133413 273668 133446 273670
rect 133510 273668 133516 273732
rect 133413 273667 133479 273668
rect 135897 273596 135963 273597
rect 138473 273596 138539 273597
rect 140865 273596 140931 273597
rect 143533 273596 143599 273597
rect 135888 273532 135894 273596
rect 135958 273594 135964 273596
rect 138472 273594 138478 273596
rect 135958 273534 136050 273594
rect 138386 273534 138478 273594
rect 135958 273532 135964 273534
rect 138472 273532 138478 273534
rect 138542 273532 138548 273596
rect 140865 273594 140926 273596
rect 140834 273592 140926 273594
rect 140834 273536 140870 273592
rect 140834 273534 140926 273536
rect 140865 273532 140926 273534
rect 140990 273532 140996 273596
rect 143504 273532 143510 273596
rect 143574 273594 143599 273596
rect 145925 273596 145991 273597
rect 266353 273596 266419 273597
rect 269757 273596 269823 273597
rect 271137 273596 271203 273597
rect 283465 273596 283531 273597
rect 421097 273596 421163 273597
rect 422845 273596 422911 273597
rect 427629 273596 427695 273597
rect 145925 273594 145958 273596
rect 143574 273592 143666 273594
rect 143594 273536 143666 273592
rect 143574 273534 143666 273536
rect 145866 273592 145958 273594
rect 145866 273536 145930 273592
rect 145866 273534 145958 273536
rect 143574 273532 143599 273534
rect 135897 273531 135963 273532
rect 138473 273531 138539 273532
rect 140865 273531 140931 273532
rect 143533 273531 143599 273532
rect 145925 273532 145958 273534
rect 146022 273532 146028 273596
rect 266353 273594 266382 273596
rect 266290 273592 266382 273594
rect 266290 273536 266358 273592
rect 266290 273534 266382 273536
rect 266353 273532 266382 273534
rect 266446 273532 266452 273596
rect 269757 273594 269782 273596
rect 269690 273592 269782 273594
rect 269690 273536 269762 273592
rect 269690 273534 269782 273536
rect 269757 273532 269782 273534
rect 269846 273532 269852 273596
rect 271136 273594 271142 273596
rect 271050 273534 271142 273594
rect 271136 273532 271142 273534
rect 271206 273532 271212 273596
rect 283465 273594 283518 273596
rect 283426 273592 283518 273594
rect 283426 273536 283470 273592
rect 283426 273534 283518 273536
rect 283465 273532 283518 273534
rect 283582 273532 283588 273596
rect 421072 273532 421078 273596
rect 421142 273594 421163 273596
rect 422840 273594 422846 273596
rect 421142 273592 421234 273594
rect 421158 273536 421234 273592
rect 421142 273534 421234 273536
rect 422754 273534 422846 273594
rect 421142 273532 421163 273534
rect 422840 273532 422846 273534
rect 422910 273532 422916 273596
rect 427600 273532 427606 273596
rect 427670 273594 427695 273596
rect 445937 273596 446003 273597
rect 445937 273594 445966 273596
rect 427670 273592 427762 273594
rect 427690 273536 427762 273592
rect 427670 273534 427762 273536
rect 445874 273592 445966 273594
rect 445874 273536 445942 273592
rect 445874 273534 445966 273536
rect 427670 273532 427695 273534
rect 145925 273531 145991 273532
rect 266353 273531 266419 273532
rect 269757 273531 269823 273532
rect 271137 273531 271203 273532
rect 283465 273531 283531 273532
rect 421097 273531 421163 273532
rect 422845 273531 422911 273532
rect 427629 273531 427695 273532
rect 445937 273532 445966 273534
rect 446030 273532 446036 273596
rect 445937 273531 446003 273532
rect 273253 273460 273319 273461
rect 273253 273458 273300 273460
rect 273208 273456 273300 273458
rect 273208 273400 273258 273456
rect 273208 273398 273300 273400
rect 273253 273396 273300 273398
rect 273364 273396 273370 273460
rect 369761 273458 369827 273461
rect 377438 273458 377444 273460
rect 369761 273456 377444 273458
rect 369761 273400 369766 273456
rect 369822 273400 377444 273456
rect 369761 273398 377444 273400
rect 273253 273395 273319 273396
rect 369761 273395 369827 273398
rect 377438 273396 377444 273398
rect 377508 273458 377514 273460
rect 377806 273458 377812 273460
rect 377508 273398 377812 273458
rect 377508 273396 377514 273398
rect 377806 273396 377812 273398
rect 377876 273396 377882 273460
rect 378174 273396 378180 273460
rect 378244 273458 378250 273460
rect 379421 273458 379487 273461
rect 378244 273456 379487 273458
rect 378244 273400 379426 273456
rect 379482 273400 379487 273456
rect 378244 273398 379487 273400
rect 378244 273396 378250 273398
rect 379421 273395 379487 273398
rect 215334 273260 215340 273324
rect 215404 273322 215410 273324
rect 215661 273322 215727 273325
rect 215404 273320 215727 273322
rect 215404 273264 215666 273320
rect 215722 273264 215727 273320
rect 215404 273262 215727 273264
rect 215404 273260 215410 273262
rect 215661 273259 215727 273262
rect 217358 273260 217364 273324
rect 217428 273322 217434 273324
rect 250662 273322 250668 273324
rect 217428 273262 250668 273322
rect 217428 273260 217434 273262
rect 250662 273260 250668 273262
rect 250732 273260 250738 273324
rect 359406 273260 359412 273324
rect 359476 273322 359482 273324
rect 430982 273322 430988 273324
rect 359476 273262 430988 273322
rect 359476 273260 359482 273262
rect 430982 273260 430988 273262
rect 431052 273260 431058 273324
rect 76005 273188 76071 273189
rect 77109 273188 77175 273189
rect 90725 273188 90791 273189
rect 93669 273188 93735 273189
rect 76005 273186 76052 273188
rect 75960 273184 76052 273186
rect 75960 273128 76010 273184
rect 75960 273126 76052 273128
rect 76005 273124 76052 273126
rect 76116 273124 76122 273188
rect 77109 273186 77156 273188
rect 77064 273184 77156 273186
rect 77064 273128 77114 273184
rect 77064 273126 77156 273128
rect 77109 273124 77156 273126
rect 77220 273124 77226 273188
rect 90725 273186 90772 273188
rect 90680 273184 90772 273186
rect 90680 273128 90730 273184
rect 90680 273126 90772 273128
rect 90725 273124 90772 273126
rect 90836 273124 90842 273188
rect 93669 273186 93716 273188
rect 93624 273184 93716 273186
rect 93624 273128 93674 273184
rect 93624 273126 93716 273128
rect 93669 273124 93716 273126
rect 93780 273124 93786 273188
rect 94221 273186 94287 273189
rect 101806 273186 101812 273188
rect 94221 273184 101812 273186
rect 94221 273128 94226 273184
rect 94282 273128 101812 273184
rect 94221 273126 101812 273128
rect 76005 273123 76071 273124
rect 77109 273123 77175 273124
rect 90725 273123 90791 273124
rect 93669 273123 93735 273124
rect 94221 273123 94287 273126
rect 101806 273124 101812 273126
rect 101876 273124 101882 273188
rect 198038 273124 198044 273188
rect 198108 273186 198114 273188
rect 318374 273186 318380 273188
rect 198108 273126 318380 273186
rect 198108 273124 198114 273126
rect 318374 273124 318380 273126
rect 318444 273124 318450 273188
rect 359590 273124 359596 273188
rect 359660 273186 359666 273188
rect 483238 273186 483244 273188
rect 359660 273126 483244 273186
rect 359660 273124 359666 273126
rect 483238 273124 483244 273126
rect 483308 273124 483314 273188
rect 47710 272988 47716 273052
rect 47780 273050 47786 273052
rect 50153 273050 50219 273053
rect 298461 273052 298527 273053
rect 423397 273052 423463 273053
rect 425237 273052 425303 273053
rect 425973 273052 426039 273053
rect 428181 273052 428247 273053
rect 468477 273052 468543 273053
rect 97022 273050 97028 273052
rect 47780 273048 97028 273050
rect 47780 272992 50158 273048
rect 50214 272992 97028 273048
rect 47780 272990 97028 272992
rect 47780 272988 47786 272990
rect 50153 272987 50219 272990
rect 97022 272988 97028 272990
rect 97092 272988 97098 273052
rect 196750 272988 196756 273052
rect 196820 273050 196826 273052
rect 298461 273050 298508 273052
rect 196820 272990 296730 273050
rect 298416 273048 298508 273050
rect 298416 272992 298466 273048
rect 298416 272990 298508 272992
rect 196820 272988 196826 272990
rect 50245 272914 50311 272917
rect 94221 272914 94287 272917
rect 94405 272916 94471 272917
rect 95877 272916 95943 272917
rect 98453 272916 98519 272917
rect 285949 272916 286015 272917
rect 288157 272916 288223 272917
rect 290917 272916 290983 272917
rect 293309 272916 293375 272917
rect 295885 272916 295951 272917
rect 94405 272914 94452 272916
rect 50245 272912 94287 272914
rect 50245 272856 50250 272912
rect 50306 272856 94226 272912
rect 94282 272856 94287 272912
rect 50245 272854 94287 272856
rect 94360 272912 94452 272914
rect 94360 272856 94410 272912
rect 94360 272854 94452 272856
rect 50245 272851 50311 272854
rect 94221 272851 94287 272854
rect 94405 272852 94452 272854
rect 94516 272852 94522 272916
rect 95877 272914 95924 272916
rect 95832 272912 95924 272914
rect 95832 272856 95882 272912
rect 95832 272854 95924 272856
rect 95877 272852 95924 272854
rect 95988 272852 95994 272916
rect 98453 272914 98500 272916
rect 98408 272912 98500 272914
rect 98408 272856 98458 272912
rect 98408 272854 98500 272856
rect 98453 272852 98500 272854
rect 98564 272852 98570 272916
rect 285949 272914 285996 272916
rect 285904 272912 285996 272914
rect 285904 272856 285954 272912
rect 285904 272854 285996 272856
rect 285949 272852 285996 272854
rect 286060 272852 286066 272916
rect 288157 272914 288204 272916
rect 288112 272912 288204 272914
rect 288112 272856 288162 272912
rect 288112 272854 288204 272856
rect 288157 272852 288204 272854
rect 288268 272852 288274 272916
rect 290917 272914 290964 272916
rect 290872 272912 290964 272914
rect 290872 272856 290922 272912
rect 290872 272854 290964 272856
rect 290917 272852 290964 272854
rect 291028 272852 291034 272916
rect 293309 272914 293356 272916
rect 293264 272912 293356 272914
rect 293264 272856 293314 272912
rect 293264 272854 293356 272856
rect 293309 272852 293356 272854
rect 293420 272852 293426 272916
rect 295885 272914 295932 272916
rect 295840 272912 295932 272914
rect 295840 272856 295890 272912
rect 295840 272854 295932 272856
rect 295885 272852 295932 272854
rect 295996 272852 296002 272916
rect 296670 272914 296730 272990
rect 298461 272988 298508 272990
rect 298572 272988 298578 273052
rect 377806 272988 377812 273052
rect 377876 273050 377882 273052
rect 423397 273050 423444 273052
rect 377876 272990 412650 273050
rect 423352 273048 423444 273050
rect 423352 272992 423402 273048
rect 423352 272990 423444 272992
rect 377876 272988 377882 272990
rect 298461 272987 298527 272988
rect 305862 272914 305868 272916
rect 296670 272854 305868 272914
rect 305862 272852 305868 272854
rect 305932 272852 305938 272916
rect 412590 272914 412650 272990
rect 423397 272988 423444 272990
rect 423508 272988 423514 273052
rect 425237 273050 425284 273052
rect 425192 273048 425284 273050
rect 425192 272992 425242 273048
rect 425192 272990 425284 272992
rect 425237 272988 425284 272990
rect 425348 272988 425354 273052
rect 425973 273050 426020 273052
rect 425928 273048 426020 273050
rect 425928 272992 425978 273048
rect 425928 272990 426020 272992
rect 425973 272988 426020 272990
rect 426084 272988 426090 273052
rect 428181 273050 428228 273052
rect 428136 273048 428228 273050
rect 428136 272992 428186 273048
rect 428136 272990 428228 272992
rect 428181 272988 428228 272990
rect 428292 272988 428298 273052
rect 468477 273050 468524 273052
rect 468432 273048 468524 273050
rect 468432 272992 468482 273048
rect 468432 272990 468524 272992
rect 468477 272988 468524 272990
rect 468588 272988 468594 273052
rect 423397 272987 423463 272988
rect 425237 272987 425303 272988
rect 425973 272987 426039 272988
rect 428181 272987 428247 272988
rect 468477 272987 468543 272988
rect 470869 272916 470935 272917
rect 478413 272916 478479 272917
rect 423806 272914 423812 272916
rect 412590 272854 423812 272914
rect 423806 272852 423812 272854
rect 423876 272852 423882 272916
rect 470869 272914 470916 272916
rect 470824 272912 470916 272914
rect 470824 272856 470874 272912
rect 470824 272854 470916 272856
rect 470869 272852 470916 272854
rect 470980 272852 470986 272916
rect 478413 272914 478460 272916
rect 478368 272912 478460 272914
rect 478368 272856 478418 272912
rect 478368 272854 478460 272856
rect 478413 272852 478460 272854
rect 478524 272852 478530 272916
rect 94405 272851 94471 272852
rect 95877 272851 95943 272852
rect 98453 272851 98519 272852
rect 285949 272851 286015 272852
rect 288157 272851 288223 272852
rect 290917 272851 290983 272852
rect 293309 272851 293375 272852
rect 295885 272851 295951 272852
rect 470869 272851 470935 272852
rect 478413 272851 478479 272852
rect 52453 272778 52519 272781
rect 300853 272780 300919 272781
rect 303429 272780 303495 272781
rect 473445 272780 473511 272781
rect 480805 272780 480871 272781
rect 103830 272778 103836 272780
rect 52453 272776 103836 272778
rect 52453 272720 52458 272776
rect 52514 272720 103836 272776
rect 52453 272718 103836 272720
rect 52453 272715 52519 272718
rect 103830 272716 103836 272718
rect 103900 272716 103906 272780
rect 300853 272778 300900 272780
rect 300808 272776 300900 272778
rect 300808 272720 300858 272776
rect 300808 272718 300900 272720
rect 300853 272716 300900 272718
rect 300964 272716 300970 272780
rect 303429 272778 303476 272780
rect 303384 272776 303476 272778
rect 303384 272720 303434 272776
rect 303384 272718 303476 272720
rect 303429 272716 303476 272718
rect 303540 272716 303546 272780
rect 473445 272778 473492 272780
rect 473400 272776 473492 272778
rect 473400 272720 473450 272776
rect 473400 272718 473492 272720
rect 473445 272716 473492 272718
rect 473556 272716 473562 272780
rect 480805 272778 480852 272780
rect 480760 272776 480852 272778
rect 480760 272720 480810 272776
rect 480760 272718 480852 272720
rect 480805 272716 480852 272718
rect 480916 272716 480922 272780
rect 300853 272715 300919 272716
rect 303429 272715 303495 272716
rect 473445 272715 473511 272716
rect 480805 272715 480871 272716
rect 59445 272642 59511 272645
rect 310973 272644 311039 272645
rect 320909 272644 320975 272645
rect 475837 272644 475903 272645
rect 485957 272644 486023 272645
rect 117998 272642 118004 272644
rect 59445 272640 118004 272642
rect 59445 272584 59450 272640
rect 59506 272584 118004 272640
rect 59445 272582 118004 272584
rect 59445 272579 59511 272582
rect 117998 272580 118004 272582
rect 118068 272580 118074 272644
rect 310973 272642 311020 272644
rect 310928 272640 311020 272642
rect 310928 272584 310978 272640
rect 310928 272582 311020 272584
rect 310973 272580 311020 272582
rect 311084 272580 311090 272644
rect 320909 272642 320956 272644
rect 320864 272640 320956 272642
rect 320864 272584 320914 272640
rect 320864 272582 320956 272584
rect 320909 272580 320956 272582
rect 321020 272580 321026 272644
rect 475837 272642 475884 272644
rect 475792 272640 475884 272642
rect 475792 272584 475842 272640
rect 475792 272582 475884 272584
rect 475837 272580 475884 272582
rect 475948 272580 475954 272644
rect 485957 272642 486004 272644
rect 485912 272640 486004 272642
rect 485912 272584 485962 272640
rect 485912 272582 486004 272584
rect 485957 272580 486004 272582
rect 486068 272580 486074 272644
rect 310973 272579 311039 272580
rect 320909 272579 320975 272580
rect 475837 272579 475903 272580
rect 485957 272579 486023 272580
rect 46013 272506 46079 272509
rect 108614 272506 108620 272508
rect 46013 272504 108620 272506
rect 46013 272448 46018 272504
rect 46074 272448 108620 272504
rect 46013 272446 108620 272448
rect 46013 272443 46079 272446
rect 108614 272444 108620 272446
rect 108684 272444 108690 272508
rect 82997 272372 83063 272373
rect 100753 272372 100819 272373
rect 82997 272370 83044 272372
rect 82952 272368 83044 272370
rect 82952 272312 83002 272368
rect 82952 272310 83044 272312
rect 82997 272308 83044 272310
rect 83108 272308 83114 272372
rect 100702 272308 100708 272372
rect 100772 272370 100819 272372
rect 100772 272368 100864 272370
rect 100814 272312 100864 272368
rect 100772 272310 100864 272312
rect 100772 272308 100819 272310
rect 82997 272307 83063 272308
rect 100753 272307 100819 272308
rect 99373 272236 99439 272237
rect 265157 272236 265223 272237
rect 401685 272236 401751 272237
rect 415853 272236 415919 272237
rect 416037 272236 416103 272237
rect 455781 272236 455847 272237
rect 99373 272234 99420 272236
rect 99328 272232 99420 272234
rect 99328 272176 99378 272232
rect 99328 272174 99420 272176
rect 99373 272172 99420 272174
rect 99484 272172 99490 272236
rect 265157 272234 265204 272236
rect 265112 272232 265204 272234
rect 265112 272176 265162 272232
rect 265112 272174 265204 272176
rect 265157 272172 265204 272174
rect 265268 272172 265274 272236
rect 401685 272234 401732 272236
rect 401640 272232 401732 272234
rect 401640 272176 401690 272232
rect 401640 272174 401732 272176
rect 401685 272172 401732 272174
rect 401796 272172 401802 272236
rect 415853 272234 415900 272236
rect 415808 272232 415900 272234
rect 415808 272176 415858 272232
rect 415808 272174 415900 272176
rect 415853 272172 415900 272174
rect 415964 272172 415970 272236
rect 416037 272232 416084 272236
rect 416148 272234 416154 272236
rect 455781 272234 455828 272236
rect 416037 272176 416042 272232
rect 416037 272172 416084 272176
rect 416148 272174 416194 272234
rect 455736 272232 455828 272234
rect 455736 272176 455786 272232
rect 455736 272174 455828 272176
rect 416148 272172 416154 272174
rect 455781 272172 455828 272174
rect 455892 272172 455898 272236
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 99373 272171 99439 272172
rect 265157 272171 265223 272172
rect 401685 272171 401751 272172
rect 415853 272171 415919 272172
rect 416037 272171 416103 272172
rect 455781 272171 455847 272172
rect 580349 272171 580415 272174
rect 583520 272084 584960 272174
rect 51625 271828 51691 271829
rect 51574 271826 51580 271828
rect 51534 271766 51580 271826
rect 51644 271824 51691 271828
rect 51686 271768 51691 271824
rect 51574 271764 51580 271766
rect 51644 271764 51691 271768
rect 51625 271763 51691 271764
rect 53005 271826 53071 271829
rect 53230 271826 53236 271828
rect 53005 271824 53236 271826
rect 53005 271768 53010 271824
rect 53066 271768 53236 271824
rect 53005 271766 53236 271768
rect 53005 271763 53071 271766
rect 53230 271764 53236 271766
rect 53300 271764 53306 271828
rect 83958 271764 83964 271828
rect 84028 271826 84034 271828
rect 84193 271826 84259 271829
rect 84028 271824 84259 271826
rect 84028 271768 84198 271824
rect 84254 271768 84259 271824
rect 84028 271766 84259 271768
rect 84028 271764 84034 271766
rect 84193 271763 84259 271766
rect 97993 271826 98059 271829
rect 98126 271826 98132 271828
rect 97993 271824 98132 271826
rect 97993 271768 97998 271824
rect 98054 271768 98132 271824
rect 97993 271766 98132 271768
rect 97993 271763 98059 271766
rect 98126 271764 98132 271766
rect 98196 271764 98202 271828
rect 102133 271826 102199 271829
rect 102726 271826 102732 271828
rect 102133 271824 102732 271826
rect 102133 271768 102138 271824
rect 102194 271768 102732 271824
rect 102133 271766 102732 271768
rect 102133 271763 102199 271766
rect 102726 271764 102732 271766
rect 102796 271764 102802 271828
rect 104893 271826 104959 271829
rect 107469 271828 107535 271829
rect 114461 271828 114527 271829
rect 105302 271826 105308 271828
rect 104893 271824 105308 271826
rect 104893 271768 104898 271824
rect 104954 271768 105308 271824
rect 104893 271766 105308 271768
rect 104893 271763 104959 271766
rect 105302 271764 105308 271766
rect 105372 271764 105378 271828
rect 107469 271824 107516 271828
rect 107580 271826 107586 271828
rect 114461 271826 114508 271828
rect 107469 271768 107474 271824
rect 107469 271764 107516 271768
rect 107580 271766 107626 271826
rect 114416 271824 114508 271826
rect 114416 271768 114466 271824
rect 114416 271766 114508 271768
rect 107580 271764 107586 271766
rect 114461 271764 114508 271766
rect 114572 271764 114578 271828
rect 123201 271826 123267 271829
rect 123518 271826 123524 271828
rect 123201 271824 123524 271826
rect 123201 271768 123206 271824
rect 123262 271768 123524 271824
rect 123201 271766 123524 271768
rect 107469 271763 107535 271764
rect 114461 271763 114527 271764
rect 123201 271763 123267 271766
rect 123518 271764 123524 271766
rect 123588 271764 123594 271828
rect 125593 271826 125659 271829
rect 125910 271826 125916 271828
rect 125593 271824 125916 271826
rect 125593 271768 125598 271824
rect 125654 271768 125916 271824
rect 125593 271766 125916 271768
rect 125593 271763 125659 271766
rect 125910 271764 125916 271766
rect 125980 271764 125986 271828
rect 129733 271826 129799 271829
rect 130878 271826 130884 271828
rect 129733 271824 130884 271826
rect 129733 271768 129738 271824
rect 129794 271768 130884 271824
rect 129733 271766 130884 271768
rect 129733 271763 129799 271766
rect 130878 271764 130884 271766
rect 130948 271764 130954 271828
rect 150934 271764 150940 271828
rect 151004 271826 151010 271828
rect 151353 271826 151419 271829
rect 151004 271824 151419 271826
rect 151004 271768 151358 271824
rect 151414 271768 151419 271824
rect 151004 271766 151419 271768
rect 151004 271764 151010 271766
rect 151353 271763 151419 271766
rect 154062 271764 154068 271828
rect 154132 271826 154138 271828
rect 154481 271826 154547 271829
rect 154132 271824 154547 271826
rect 154132 271768 154486 271824
rect 154542 271768 154547 271824
rect 154132 271766 154547 271768
rect 154132 271764 154138 271766
rect 154481 271763 154547 271766
rect 158478 271764 158484 271828
rect 158548 271826 158554 271828
rect 158621 271826 158687 271829
rect 158548 271824 158687 271826
rect 158548 271768 158626 271824
rect 158682 271768 158687 271824
rect 158548 271766 158687 271768
rect 158548 271764 158554 271766
rect 158621 271763 158687 271766
rect 212809 271826 212875 271829
rect 213361 271826 213427 271829
rect 263593 271828 263659 271829
rect 212809 271824 213427 271826
rect 212809 271768 212814 271824
rect 212870 271768 213366 271824
rect 213422 271768 213427 271824
rect 212809 271766 213427 271768
rect 212809 271763 212875 271766
rect 213361 271763 213427 271766
rect 263542 271764 263548 271828
rect 263612 271826 263659 271828
rect 270493 271826 270559 271829
rect 270902 271826 270908 271828
rect 263612 271824 263704 271826
rect 263654 271768 263704 271824
rect 263612 271766 263704 271768
rect 270493 271824 270908 271826
rect 270493 271768 270498 271824
rect 270554 271768 270908 271824
rect 270493 271766 270908 271768
rect 263612 271764 263659 271766
rect 263593 271763 263659 271764
rect 270493 271763 270559 271766
rect 270902 271764 270908 271766
rect 270972 271764 270978 271828
rect 271873 271826 271939 271829
rect 272558 271826 272564 271828
rect 271873 271824 272564 271826
rect 271873 271768 271878 271824
rect 271934 271768 272564 271824
rect 271873 271766 272564 271768
rect 271873 271763 271939 271766
rect 272558 271764 272564 271766
rect 272628 271764 272634 271828
rect 276013 271826 276079 271829
rect 276974 271826 276980 271828
rect 276013 271824 276980 271826
rect 276013 271768 276018 271824
rect 276074 271768 276980 271824
rect 276013 271766 276980 271768
rect 276013 271763 276079 271766
rect 276974 271764 276980 271766
rect 277044 271764 277050 271828
rect 277945 271826 278011 271829
rect 278446 271826 278452 271828
rect 277945 271824 278452 271826
rect 277945 271768 277950 271824
rect 278006 271768 278452 271824
rect 277945 271766 278452 271768
rect 277945 271763 278011 271766
rect 278446 271764 278452 271766
rect 278516 271764 278522 271828
rect 280153 271826 280219 271829
rect 280838 271826 280844 271828
rect 280153 271824 280844 271826
rect 280153 271768 280158 271824
rect 280214 271768 280844 271824
rect 280153 271766 280844 271768
rect 280153 271763 280219 271766
rect 280838 271764 280844 271766
rect 280908 271764 280914 271828
rect 307753 271826 307819 271829
rect 308622 271826 308628 271828
rect 307753 271824 308628 271826
rect 307753 271768 307758 271824
rect 307814 271768 308628 271824
rect 307753 271766 308628 271768
rect 307753 271763 307819 271766
rect 308622 271764 308628 271766
rect 308692 271764 308698 271828
rect 343398 271764 343404 271828
rect 343468 271826 343474 271828
rect 343541 271826 343607 271829
rect 343468 271824 343607 271826
rect 343468 271768 343546 271824
rect 343602 271768 343607 271824
rect 343468 271766 343607 271768
rect 343468 271764 343474 271766
rect 343541 271763 343607 271766
rect 427813 271826 427879 271829
rect 428590 271826 428596 271828
rect 427813 271824 428596 271826
rect 427813 271768 427818 271824
rect 427874 271768 428596 271824
rect 427813 271766 428596 271768
rect 427813 271763 427879 271766
rect 428590 271764 428596 271766
rect 428660 271764 428666 271828
rect 430573 271826 430639 271829
rect 431166 271826 431172 271828
rect 430573 271824 431172 271826
rect 430573 271768 430578 271824
rect 430634 271768 431172 271824
rect 430573 271766 431172 271768
rect 430573 271763 430639 271766
rect 431166 271764 431172 271766
rect 431236 271764 431242 271828
rect 432045 271826 432111 271829
rect 433333 271828 433399 271829
rect 432270 271826 432276 271828
rect 432045 271824 432276 271826
rect 432045 271768 432050 271824
rect 432106 271768 432276 271824
rect 432045 271766 432276 271768
rect 432045 271763 432111 271766
rect 432270 271764 432276 271766
rect 432340 271764 432346 271828
rect 433333 271826 433380 271828
rect 433288 271824 433380 271826
rect 433288 271768 433338 271824
rect 433288 271766 433380 271768
rect 433333 271764 433380 271766
rect 433444 271764 433450 271828
rect 434713 271826 434779 271829
rect 435950 271826 435956 271828
rect 434713 271824 435956 271826
rect 434713 271768 434718 271824
rect 434774 271768 435956 271824
rect 434713 271766 435956 271768
rect 433333 271763 433399 271764
rect 434713 271763 434779 271766
rect 435950 271764 435956 271766
rect 436020 271764 436026 271828
rect 437473 271826 437539 271829
rect 438526 271826 438532 271828
rect 437473 271824 438532 271826
rect 437473 271768 437478 271824
rect 437534 271768 438532 271824
rect 437473 271766 438532 271768
rect 437473 271763 437539 271766
rect 438526 271764 438532 271766
rect 438596 271764 438602 271828
rect 442993 271826 443059 271829
rect 443494 271826 443500 271828
rect 442993 271824 443500 271826
rect 442993 271768 442998 271824
rect 443054 271768 443500 271824
rect 442993 271766 443500 271768
rect 442993 271763 443059 271766
rect 443494 271764 443500 271766
rect 443564 271764 443570 271828
rect 447133 271826 447199 271829
rect 448278 271826 448284 271828
rect 447133 271824 448284 271826
rect 447133 271768 447138 271824
rect 447194 271768 448284 271824
rect 447133 271766 448284 271768
rect 447133 271763 447199 271766
rect 448278 271764 448284 271766
rect 448348 271764 448354 271828
rect 449893 271826 449959 271829
rect 451038 271826 451044 271828
rect 449893 271824 451044 271826
rect 449893 271768 449898 271824
rect 449954 271768 451044 271824
rect 449893 271766 451044 271768
rect 449893 271763 449959 271766
rect 451038 271764 451044 271766
rect 451108 271764 451114 271828
rect 452653 271826 452719 271829
rect 453430 271826 453436 271828
rect 452653 271824 453436 271826
rect 452653 271768 452658 271824
rect 452714 271768 453436 271824
rect 452653 271766 453436 271768
rect 452653 271763 452719 271766
rect 453430 271764 453436 271766
rect 453500 271764 453506 271828
rect 458173 271826 458239 271829
rect 458398 271826 458404 271828
rect 458173 271824 458404 271826
rect 458173 271768 458178 271824
rect 458234 271768 458404 271824
rect 458173 271766 458404 271768
rect 458173 271763 458239 271766
rect 458398 271764 458404 271766
rect 458468 271764 458474 271828
rect 49049 271690 49115 271693
rect 81934 271690 81940 271692
rect 49049 271688 81940 271690
rect 49049 271632 49054 271688
rect 49110 271632 81940 271688
rect 49049 271630 81940 271632
rect 49049 271627 49115 271630
rect 81934 271628 81940 271630
rect 82004 271628 82010 271692
rect 100753 271690 100819 271693
rect 101070 271690 101076 271692
rect 100753 271688 101076 271690
rect 100753 271632 100758 271688
rect 100814 271632 101076 271688
rect 100753 271630 101076 271632
rect 100753 271627 100819 271630
rect 101070 271628 101076 271630
rect 101140 271628 101146 271692
rect 110413 271690 110479 271693
rect 111006 271690 111012 271692
rect 110413 271688 111012 271690
rect 110413 271632 110418 271688
rect 110474 271632 111012 271688
rect 110413 271630 111012 271632
rect 110413 271627 110479 271630
rect 111006 271628 111012 271630
rect 111076 271628 111082 271692
rect 120073 271690 120139 271693
rect 120758 271690 120764 271692
rect 120073 271688 120764 271690
rect 120073 271632 120078 271688
rect 120134 271632 120764 271688
rect 120073 271630 120764 271632
rect 120073 271627 120139 271630
rect 120758 271628 120764 271630
rect 120828 271628 120834 271692
rect 128353 271690 128419 271693
rect 128670 271690 128676 271692
rect 128353 271688 128676 271690
rect 128353 271632 128358 271688
rect 128414 271632 128676 271688
rect 128353 271630 128676 271632
rect 128353 271627 128419 271630
rect 128670 271628 128676 271630
rect 128740 271628 128746 271692
rect 155902 271628 155908 271692
rect 155972 271690 155978 271692
rect 157241 271690 157307 271693
rect 155972 271688 157307 271690
rect 155972 271632 157246 271688
rect 157302 271632 157307 271688
rect 155972 271630 157307 271632
rect 155972 271628 155978 271630
rect 157241 271627 157307 271630
rect 160870 271628 160876 271692
rect 160940 271690 160946 271692
rect 161289 271690 161355 271693
rect 160940 271688 161355 271690
rect 160940 271632 161294 271688
rect 161350 271632 161355 271688
rect 160940 271630 161355 271632
rect 160940 271628 160946 271630
rect 161289 271627 161355 271630
rect 163446 271628 163452 271692
rect 163516 271690 163522 271692
rect 164141 271690 164207 271693
rect 163516 271688 164207 271690
rect 163516 271632 164146 271688
rect 164202 271632 164207 271688
rect 163516 271630 164207 271632
rect 163516 271628 163522 271630
rect 164141 271627 164207 271630
rect 166022 271628 166028 271692
rect 166092 271690 166098 271692
rect 166901 271690 166967 271693
rect 166092 271688 166967 271690
rect 166092 271632 166906 271688
rect 166962 271632 166967 271688
rect 166092 271630 166967 271632
rect 166092 271628 166098 271630
rect 166901 271627 166967 271630
rect 183134 271628 183140 271692
rect 183204 271690 183210 271692
rect 183461 271690 183527 271693
rect 183204 271688 183527 271690
rect 183204 271632 183466 271688
rect 183522 271632 183527 271688
rect 183204 271630 183527 271632
rect 183204 271628 183210 271630
rect 183461 271627 183527 271630
rect 212073 271690 212139 271693
rect 315062 271690 315068 271692
rect 212073 271688 315068 271690
rect 212073 271632 212078 271688
rect 212134 271632 315068 271688
rect 212073 271630 315068 271632
rect 212073 271627 212139 271630
rect 315062 271628 315068 271630
rect 315132 271628 315138 271692
rect 379053 271690 379119 271693
rect 465942 271690 465948 271692
rect 379053 271688 465948 271690
rect 379053 271632 379058 271688
rect 379114 271632 465948 271688
rect 379053 271630 465948 271632
rect 379053 271627 379119 271630
rect 465942 271628 465948 271630
rect 466012 271628 466018 271692
rect 503110 271628 503116 271692
rect 503180 271690 503186 271692
rect 503621 271690 503687 271693
rect 503180 271688 503687 271690
rect 503180 271632 503626 271688
rect 503682 271632 503687 271688
rect 503180 271630 503687 271632
rect 503180 271628 503186 271630
rect 503621 271627 503687 271630
rect 47669 271554 47735 271557
rect 115933 271556 115999 271557
rect 79542 271554 79548 271556
rect 47669 271552 79548 271554
rect 47669 271496 47674 271552
rect 47730 271496 79548 271552
rect 47669 271494 79548 271496
rect 47669 271491 47735 271494
rect 79542 271492 79548 271494
rect 79612 271492 79618 271556
rect 115933 271554 115980 271556
rect 115888 271552 115980 271554
rect 115888 271496 115938 271552
rect 115888 271494 115980 271496
rect 115933 271492 115980 271494
rect 116044 271492 116050 271556
rect 117313 271554 117379 271557
rect 118366 271554 118372 271556
rect 117313 271552 118372 271554
rect 117313 271496 117318 271552
rect 117374 271496 118372 271552
rect 117313 271494 118372 271496
rect 115933 271491 115999 271492
rect 117313 271491 117379 271494
rect 118366 271492 118372 271494
rect 118436 271492 118442 271556
rect 217174 271492 217180 271556
rect 217244 271554 217250 271556
rect 273478 271554 273484 271556
rect 217244 271494 273484 271554
rect 217244 271492 217250 271494
rect 273478 271492 273484 271494
rect 273548 271492 273554 271556
rect 276013 271554 276079 271557
rect 276238 271554 276244 271556
rect 276013 271552 276244 271554
rect 276013 271496 276018 271552
rect 276074 271496 276244 271552
rect 276013 271494 276244 271496
rect 276013 271491 276079 271494
rect 276238 271492 276244 271494
rect 276308 271492 276314 271556
rect 376293 271554 376359 271557
rect 460974 271554 460980 271556
rect 376293 271552 460980 271554
rect 376293 271496 376298 271552
rect 376354 271496 460980 271552
rect 376293 271494 460980 271496
rect 376293 271491 376359 271494
rect 460974 271492 460980 271494
rect 461044 271492 461050 271556
rect 47853 271418 47919 271421
rect 78254 271418 78260 271420
rect 47853 271416 78260 271418
rect 47853 271360 47858 271416
rect 47914 271360 78260 271416
rect 47853 271358 78260 271360
rect 47853 271355 47919 271358
rect 78254 271356 78260 271358
rect 78324 271356 78330 271420
rect 103513 271418 103579 271421
rect 113173 271420 113239 271421
rect 103830 271418 103836 271420
rect 103513 271416 103836 271418
rect 103513 271360 103518 271416
rect 103574 271360 103836 271416
rect 103513 271358 103836 271360
rect 103513 271355 103579 271358
rect 103830 271356 103836 271358
rect 103900 271356 103906 271420
rect 113173 271416 113220 271420
rect 113284 271418 113290 271420
rect 213361 271418 213427 271421
rect 236494 271418 236500 271420
rect 113173 271360 113178 271416
rect 113173 271356 113220 271360
rect 113284 271358 113330 271418
rect 213361 271416 236500 271418
rect 213361 271360 213366 271416
rect 213422 271360 236500 271416
rect 213361 271358 236500 271360
rect 113284 271356 113290 271358
rect 113173 271355 113239 271356
rect 213361 271355 213427 271358
rect 236494 271356 236500 271358
rect 236564 271356 236570 271420
rect 260833 271418 260899 271421
rect 260966 271418 260972 271420
rect 260833 271416 260972 271418
rect 260833 271360 260838 271416
rect 260894 271360 260972 271416
rect 260833 271358 260972 271360
rect 260833 271355 260899 271358
rect 260966 271356 260972 271358
rect 261036 271356 261042 271420
rect 267825 271418 267891 271421
rect 268326 271418 268332 271420
rect 267825 271416 268332 271418
rect 267825 271360 267830 271416
rect 267886 271360 268332 271416
rect 267825 271358 268332 271360
rect 267825 271355 267891 271358
rect 268326 271356 268332 271358
rect 268396 271356 268402 271420
rect 343214 271356 343220 271420
rect 343284 271418 343290 271420
rect 343541 271418 343607 271421
rect 343284 271416 343607 271418
rect 343284 271360 343546 271416
rect 343602 271360 343607 271416
rect 343284 271358 343607 271360
rect 343284 271356 343290 271358
rect 343541 271355 343607 271358
rect 377254 271356 377260 271420
rect 377324 271418 377330 271420
rect 408166 271418 408172 271420
rect 377324 271358 408172 271418
rect 377324 271356 377330 271358
rect 408166 271356 408172 271358
rect 408236 271356 408242 271420
rect 433333 271418 433399 271421
rect 433558 271418 433564 271420
rect 433333 271416 433564 271418
rect 433333 271360 433338 271416
rect 433394 271360 433564 271416
rect 433333 271358 433564 271360
rect 433333 271355 433399 271358
rect 433558 271356 433564 271358
rect 433628 271356 433634 271420
rect 440233 271418 440299 271421
rect 440918 271418 440924 271420
rect 440233 271416 440924 271418
rect 440233 271360 440238 271416
rect 440294 271360 440924 271416
rect 440233 271358 440924 271360
rect 440233 271355 440299 271358
rect 440918 271356 440924 271358
rect 440988 271356 440994 271420
rect 104893 271282 104959 271285
rect 105854 271282 105860 271284
rect 104893 271280 105860 271282
rect 104893 271224 104898 271280
rect 104954 271224 105860 271280
rect 104893 271222 105860 271224
rect 104893 271219 104959 271222
rect 105854 271220 105860 271222
rect 105924 271220 105930 271284
rect 107653 271282 107719 271285
rect 108246 271282 108252 271284
rect 107653 271280 108252 271282
rect 107653 271224 107658 271280
rect 107714 271224 108252 271280
rect 107653 271222 108252 271224
rect 107653 271219 107719 271222
rect 108246 271220 108252 271222
rect 108316 271220 108322 271284
rect 118693 271282 118759 271285
rect 119102 271282 119108 271284
rect 118693 271280 119108 271282
rect 118693 271224 118698 271280
rect 118754 271224 119108 271280
rect 118693 271222 119108 271224
rect 118693 271219 118759 271222
rect 119102 271220 119108 271222
rect 119172 271220 119178 271284
rect 258257 271282 258323 271285
rect 258390 271282 258396 271284
rect 258257 271280 258396 271282
rect 258257 271224 258262 271280
rect 258318 271224 258396 271280
rect 258257 271222 258396 271224
rect 258257 271219 258323 271222
rect 258390 271220 258396 271222
rect 258460 271220 258466 271284
rect 264973 271282 265039 271285
rect 265934 271282 265940 271284
rect 264973 271280 265940 271282
rect 264973 271224 264978 271280
rect 265034 271224 265940 271280
rect 264973 271222 265940 271224
rect 264973 271219 265039 271222
rect 265934 271220 265940 271222
rect 266004 271220 266010 271284
rect 275318 271220 275324 271284
rect 275388 271282 275394 271284
rect 275921 271282 275987 271285
rect 275388 271280 275987 271282
rect 275388 271224 275926 271280
rect 275982 271224 275987 271280
rect 275388 271222 275987 271224
rect 275388 271220 275394 271222
rect 275921 271219 275987 271222
rect 278078 271220 278084 271284
rect 278148 271282 278154 271284
rect 278681 271282 278747 271285
rect 278148 271280 278747 271282
rect 278148 271224 278686 271280
rect 278742 271224 278747 271280
rect 278148 271222 278747 271224
rect 278148 271220 278154 271222
rect 278681 271219 278747 271222
rect 374361 271282 374427 271285
rect 396022 271282 396028 271284
rect 374361 271280 396028 271282
rect 374361 271224 374366 271280
rect 374422 271224 396028 271280
rect 374361 271222 396028 271224
rect 374361 271219 374427 271222
rect 396022 271220 396028 271222
rect 396092 271220 396098 271284
rect 439262 271220 439268 271284
rect 439332 271282 439338 271284
rect 440141 271282 440207 271285
rect 439332 271280 440207 271282
rect 439332 271224 440146 271280
rect 440202 271224 440207 271280
rect 439332 271222 440207 271224
rect 439332 271220 439338 271222
rect 440141 271219 440207 271222
rect 503478 271220 503484 271284
rect 503548 271282 503554 271284
rect 503621 271282 503687 271285
rect 503548 271280 503687 271282
rect 503548 271224 503626 271280
rect 503682 271224 503687 271280
rect 503548 271222 503687 271224
rect 503548 271220 503554 271222
rect 503621 271219 503687 271222
rect 53833 271146 53899 271149
rect 54385 271146 54451 271149
rect 62113 271146 62179 271149
rect 53833 271144 62179 271146
rect 53833 271088 53838 271144
rect 53894 271088 54390 271144
rect 54446 271088 62118 271144
rect 62174 271088 62179 271144
rect 53833 271086 62179 271088
rect 53833 271083 53899 271086
rect 54385 271083 54451 271086
rect 62113 271083 62179 271086
rect 111793 271146 111859 271149
rect 112110 271146 112116 271148
rect 111793 271144 112116 271146
rect 111793 271088 111798 271144
rect 111854 271088 112116 271144
rect 111793 271086 112116 271088
rect 111793 271083 111859 271086
rect 112110 271084 112116 271086
rect 112180 271084 112186 271148
rect 247033 271146 247099 271149
rect 248270 271146 248276 271148
rect 247033 271144 248276 271146
rect 247033 271088 247038 271144
rect 247094 271088 248276 271144
rect 247033 271086 248276 271088
rect 247033 271083 247099 271086
rect 248270 271084 248276 271086
rect 248340 271084 248346 271148
rect 252553 271146 252619 271149
rect 253606 271146 253612 271148
rect 252553 271144 253612 271146
rect 252553 271088 252558 271144
rect 252614 271088 253612 271144
rect 252553 271086 253612 271088
rect 252553 271083 252619 271086
rect 253606 271084 253612 271086
rect 253676 271084 253682 271148
rect 255313 271146 255379 271149
rect 256182 271146 256188 271148
rect 255313 271144 256188 271146
rect 255313 271088 255318 271144
rect 255374 271088 256188 271144
rect 255313 271086 256188 271088
rect 255313 271083 255379 271086
rect 256182 271084 256188 271086
rect 256252 271084 256258 271148
rect 313273 271146 313339 271149
rect 313406 271146 313412 271148
rect 313273 271144 313412 271146
rect 313273 271088 313278 271144
rect 313334 271088 313412 271144
rect 313273 271086 313412 271088
rect 313273 271083 313339 271086
rect 313406 271084 313412 271086
rect 313476 271084 313482 271148
rect 379789 271146 379855 271149
rect 397126 271146 397132 271148
rect 379789 271144 397132 271146
rect 379789 271088 379794 271144
rect 379850 271088 397132 271144
rect 379789 271086 397132 271088
rect 379789 271083 379855 271086
rect 397126 271084 397132 271086
rect 397196 271084 397202 271148
rect 409873 271146 409939 271149
rect 410742 271146 410748 271148
rect 409873 271144 410748 271146
rect 409873 271088 409878 271144
rect 409934 271088 410748 271144
rect 409873 271086 410748 271088
rect 409873 271083 409939 271086
rect 410742 271084 410748 271086
rect 410812 271084 410818 271148
rect 412725 271146 412791 271149
rect 413686 271146 413692 271148
rect 412725 271144 413692 271146
rect 412725 271088 412730 271144
rect 412786 271088 413692 271144
rect 412725 271086 413692 271088
rect 412725 271083 412791 271086
rect 413686 271084 413692 271086
rect 413756 271084 413762 271148
rect 418153 271146 418219 271149
rect 418470 271146 418476 271148
rect 418153 271144 418476 271146
rect 418153 271088 418158 271144
rect 418214 271088 418476 271144
rect 418153 271086 418476 271088
rect 418153 271083 418219 271086
rect 418470 271084 418476 271086
rect 418540 271084 418546 271148
rect 46565 271010 46631 271013
rect 88333 271012 88399 271013
rect 80462 271010 80468 271012
rect 46565 271008 80468 271010
rect 46565 270952 46570 271008
rect 46626 270952 80468 271008
rect 46565 270950 80468 270952
rect 46565 270947 46631 270950
rect 80462 270948 80468 270950
rect 80532 270948 80538 271012
rect 88333 271010 88380 271012
rect 88288 271008 88380 271010
rect 88288 270952 88338 271008
rect 88288 270950 88380 270952
rect 88333 270948 88380 270950
rect 88444 270948 88450 271012
rect 89713 271010 89779 271013
rect 90030 271010 90036 271012
rect 89713 271008 90036 271010
rect 89713 270952 89718 271008
rect 89774 270952 90036 271008
rect 89713 270950 90036 270952
rect 88333 270947 88399 270948
rect 89713 270947 89779 270950
rect 90030 270948 90036 270950
rect 90100 270948 90106 271012
rect 114553 271010 114619 271013
rect 115790 271010 115796 271012
rect 114553 271008 115796 271010
rect 114553 270952 114558 271008
rect 114614 270952 115796 271008
rect 114553 270950 115796 270952
rect 114553 270947 114619 270950
rect 115790 270948 115796 270950
rect 115860 270948 115866 271012
rect 207749 271010 207815 271013
rect 325550 271010 325556 271012
rect 207749 271008 325556 271010
rect 207749 270952 207754 271008
rect 207810 270952 325556 271008
rect 207749 270950 325556 270952
rect 207749 270947 207815 270950
rect 325550 270948 325556 270950
rect 325620 270948 325626 271012
rect 373533 271010 373599 271013
rect 462630 271010 462636 271012
rect 373533 271008 462636 271010
rect 373533 270952 373538 271008
rect 373594 270952 462636 271008
rect 373533 270950 462636 270952
rect 373533 270947 373599 270950
rect 462630 270948 462636 270950
rect 462700 270948 462706 271012
rect 85573 270874 85639 270877
rect 86534 270874 86540 270876
rect 85573 270872 86540 270874
rect 85573 270816 85578 270872
rect 85634 270816 86540 270872
rect 85573 270814 86540 270816
rect 85573 270811 85639 270814
rect 86534 270812 86540 270814
rect 86604 270812 86610 270876
rect 88333 270874 88399 270877
rect 88742 270874 88748 270876
rect 88333 270872 88748 270874
rect 88333 270816 88338 270872
rect 88394 270816 88748 270872
rect 88333 270814 88748 270816
rect 88333 270811 88399 270814
rect 88742 270812 88748 270814
rect 88812 270812 88818 270876
rect 92473 270874 92539 270877
rect 93342 270874 93348 270876
rect 92473 270872 93348 270874
rect 92473 270816 92478 270872
rect 92534 270816 93348 270872
rect 92473 270814 93348 270816
rect 92473 270811 92539 270814
rect 93342 270812 93348 270814
rect 93412 270812 93418 270876
rect 106273 270874 106339 270877
rect 106406 270874 106412 270876
rect 106273 270872 106412 270874
rect 106273 270816 106278 270872
rect 106334 270816 106412 270872
rect 106273 270814 106412 270816
rect 106273 270811 106339 270814
rect 106406 270812 106412 270814
rect 106476 270812 106482 270876
rect 115933 270874 115999 270877
rect 116894 270874 116900 270876
rect 115933 270872 116900 270874
rect 115933 270816 115938 270872
rect 115994 270816 116900 270872
rect 115933 270814 116900 270816
rect 115933 270811 115999 270814
rect 116894 270812 116900 270814
rect 116964 270812 116970 270876
rect 147673 270874 147739 270877
rect 148542 270874 148548 270876
rect 147673 270872 148548 270874
rect 147673 270816 147678 270872
rect 147734 270816 148548 270872
rect 147673 270814 148548 270816
rect 147673 270811 147739 270814
rect 148542 270812 148548 270814
rect 148612 270812 148618 270876
rect 253933 270874 253999 270877
rect 254526 270874 254532 270876
rect 253933 270872 254532 270874
rect 253933 270816 253938 270872
rect 253994 270816 254532 270872
rect 253933 270814 254532 270816
rect 253933 270811 253999 270814
rect 254526 270812 254532 270814
rect 254596 270812 254602 270876
rect 278998 270812 279004 270876
rect 279068 270874 279074 270876
rect 280061 270874 280127 270877
rect 279068 270872 280127 270874
rect 279068 270816 280066 270872
rect 280122 270816 280127 270872
rect 279068 270814 280127 270816
rect 279068 270812 279074 270814
rect 280061 270811 280127 270814
rect 405733 270874 405799 270877
rect 434713 270876 434779 270877
rect 406510 270874 406516 270876
rect 405733 270872 406516 270874
rect 405733 270816 405738 270872
rect 405794 270816 406516 270872
rect 405733 270814 406516 270816
rect 405733 270811 405799 270814
rect 406510 270812 406516 270814
rect 406580 270812 406586 270876
rect 434662 270812 434668 270876
rect 434732 270874 434779 270876
rect 436093 270874 436159 270877
rect 436870 270874 436876 270876
rect 434732 270872 434824 270874
rect 434774 270816 434824 270872
rect 434732 270814 434824 270816
rect 436093 270872 436876 270874
rect 436093 270816 436098 270872
rect 436154 270816 436876 270872
rect 436093 270814 436876 270816
rect 434732 270812 434779 270814
rect 434713 270811 434779 270812
rect 436093 270811 436159 270814
rect 436870 270812 436876 270814
rect 436940 270812 436946 270876
rect 437473 270874 437539 270877
rect 438342 270874 438348 270876
rect 437473 270872 438348 270874
rect 437473 270816 437478 270872
rect 437534 270816 438348 270872
rect 437473 270814 438348 270816
rect 437473 270811 437539 270814
rect 438342 270812 438348 270814
rect 438412 270812 438418 270876
rect 244222 270676 244228 270740
rect 244292 270738 244298 270740
rect 244365 270738 244431 270741
rect 251265 270740 251331 270741
rect 244292 270736 244431 270738
rect 244292 270680 244370 270736
rect 244426 270680 244431 270736
rect 244292 270678 244431 270680
rect 244292 270676 244298 270678
rect 244365 270675 244431 270678
rect 251214 270676 251220 270740
rect 251284 270738 251331 270740
rect 255313 270738 255379 270741
rect 255814 270738 255820 270740
rect 251284 270736 251376 270738
rect 251326 270680 251376 270736
rect 251284 270678 251376 270680
rect 255313 270736 255820 270738
rect 255313 270680 255318 270736
rect 255374 270680 255820 270736
rect 255313 270678 255820 270680
rect 251284 270676 251331 270678
rect 251265 270675 251331 270676
rect 255313 270675 255379 270678
rect 255814 270676 255820 270678
rect 255884 270676 255890 270740
rect 259545 270738 259611 270741
rect 411345 270740 411411 270741
rect 260598 270738 260604 270740
rect 259545 270736 260604 270738
rect 259545 270680 259550 270736
rect 259606 270680 260604 270736
rect 259545 270678 260604 270680
rect 259545 270675 259611 270678
rect 260598 270676 260604 270678
rect 260668 270676 260674 270740
rect 411294 270676 411300 270740
rect 411364 270738 411411 270740
rect 429193 270738 429259 270741
rect 429694 270738 429700 270740
rect 411364 270736 411456 270738
rect 411406 270680 411456 270736
rect 411364 270678 411456 270680
rect 429193 270736 429700 270738
rect 429193 270680 429198 270736
rect 429254 270680 429700 270736
rect 429193 270678 429700 270680
rect 411364 270676 411411 270678
rect 411345 270675 411411 270676
rect 429193 270675 429259 270678
rect 429694 270676 429700 270678
rect 429764 270676 429770 270740
rect 434805 270738 434871 270741
rect 435766 270738 435772 270740
rect 434805 270736 435772 270738
rect 434805 270680 434810 270736
rect 434866 270680 435772 270736
rect 434805 270678 435772 270680
rect 434805 270675 434871 270678
rect 435766 270676 435772 270678
rect 435836 270676 435842 270740
rect 84653 270604 84719 270605
rect 84653 270602 84700 270604
rect 84608 270600 84700 270602
rect 84608 270544 84658 270600
rect 84608 270542 84700 270544
rect 84653 270540 84700 270542
rect 84764 270540 84770 270604
rect 86953 270602 87019 270605
rect 87638 270602 87644 270604
rect 86953 270600 87644 270602
rect 86953 270544 86958 270600
rect 87014 270544 87644 270600
rect 86953 270542 87644 270544
rect 84653 270539 84719 270540
rect 86953 270539 87019 270542
rect 87638 270540 87644 270542
rect 87708 270540 87714 270604
rect 91093 270602 91159 270605
rect 91318 270602 91324 270604
rect 91093 270600 91324 270602
rect 91093 270544 91098 270600
rect 91154 270544 91324 270600
rect 91093 270542 91324 270544
rect 91093 270539 91159 270542
rect 91318 270540 91324 270542
rect 91388 270540 91394 270604
rect 109033 270602 109099 270605
rect 109534 270602 109540 270604
rect 109033 270600 109540 270602
rect 109033 270544 109038 270600
rect 109094 270544 109540 270600
rect 109033 270542 109540 270544
rect 109033 270539 109099 270542
rect 109534 270540 109540 270542
rect 109604 270540 109610 270604
rect 110413 270602 110479 270605
rect 183461 270604 183527 270605
rect 111190 270602 111196 270604
rect 110413 270600 111196 270602
rect 110413 270544 110418 270600
rect 110474 270544 111196 270600
rect 110413 270542 111196 270544
rect 110413 270539 110479 270542
rect 111190 270540 111196 270542
rect 111260 270540 111266 270604
rect 183461 270602 183508 270604
rect 183416 270600 183508 270602
rect 183416 270544 183466 270600
rect 183416 270542 183508 270544
rect 183461 270540 183508 270542
rect 183572 270540 183578 270604
rect 235993 270602 236059 270605
rect 237046 270602 237052 270604
rect 235993 270600 237052 270602
rect 235993 270544 235998 270600
rect 236054 270544 237052 270600
rect 235993 270542 237052 270544
rect 183461 270539 183527 270540
rect 235993 270539 236059 270542
rect 237046 270540 237052 270542
rect 237116 270540 237122 270604
rect 237373 270602 237439 270605
rect 242893 270604 242959 270605
rect 238150 270602 238156 270604
rect 237373 270600 238156 270602
rect 237373 270544 237378 270600
rect 237434 270544 238156 270600
rect 237373 270542 238156 270544
rect 237373 270539 237439 270542
rect 238150 270540 238156 270542
rect 238220 270540 238226 270604
rect 242893 270602 242940 270604
rect 242848 270600 242940 270602
rect 242848 270544 242898 270600
rect 242848 270542 242940 270544
rect 242893 270540 242940 270542
rect 243004 270540 243010 270604
rect 244273 270602 244339 270605
rect 245326 270602 245332 270604
rect 244273 270600 245332 270602
rect 244273 270544 244278 270600
rect 244334 270544 245332 270600
rect 244273 270542 245332 270544
rect 242893 270539 242959 270540
rect 244273 270539 244339 270542
rect 245326 270540 245332 270542
rect 245396 270540 245402 270604
rect 245653 270602 245719 270605
rect 246430 270602 246436 270604
rect 245653 270600 246436 270602
rect 245653 270544 245658 270600
rect 245714 270544 246436 270600
rect 245653 270542 246436 270544
rect 245653 270539 245719 270542
rect 246430 270540 246436 270542
rect 246500 270540 246506 270604
rect 247033 270602 247099 270605
rect 247718 270602 247724 270604
rect 247033 270600 247724 270602
rect 247033 270544 247038 270600
rect 247094 270544 247724 270600
rect 247033 270542 247724 270544
rect 247033 270539 247099 270542
rect 247718 270540 247724 270542
rect 247788 270540 247794 270604
rect 248505 270602 248571 270605
rect 248638 270602 248644 270604
rect 248505 270600 248644 270602
rect 248505 270544 248510 270600
rect 248566 270544 248644 270600
rect 248505 270542 248644 270544
rect 248505 270539 248571 270542
rect 248638 270540 248644 270542
rect 248708 270540 248714 270604
rect 249793 270602 249859 270605
rect 250110 270602 250116 270604
rect 249793 270600 250116 270602
rect 249793 270544 249798 270600
rect 249854 270544 250116 270600
rect 249793 270542 250116 270544
rect 249793 270539 249859 270542
rect 250110 270540 250116 270542
rect 250180 270540 250186 270604
rect 251173 270602 251239 270605
rect 252318 270602 252324 270604
rect 251173 270600 252324 270602
rect 251173 270544 251178 270600
rect 251234 270544 252324 270600
rect 251173 270542 252324 270544
rect 251173 270539 251239 270542
rect 252318 270540 252324 270542
rect 252388 270540 252394 270604
rect 252553 270602 252619 270605
rect 253422 270602 253428 270604
rect 252553 270600 253428 270602
rect 252553 270544 252558 270600
rect 252614 270544 253428 270600
rect 252553 270542 253428 270544
rect 252553 270539 252619 270542
rect 253422 270540 253428 270542
rect 253492 270540 253498 270604
rect 256693 270602 256759 270605
rect 256918 270602 256924 270604
rect 256693 270600 256924 270602
rect 256693 270544 256698 270600
rect 256754 270544 256924 270600
rect 256693 270542 256924 270544
rect 256693 270539 256759 270542
rect 256918 270540 256924 270542
rect 256988 270540 256994 270604
rect 258073 270602 258139 270605
rect 259453 270604 259519 270605
rect 258390 270602 258396 270604
rect 258073 270600 258396 270602
rect 258073 270544 258078 270600
rect 258134 270544 258396 270600
rect 258073 270542 258396 270544
rect 258073 270539 258139 270542
rect 258390 270540 258396 270542
rect 258460 270540 258466 270604
rect 259453 270602 259500 270604
rect 259408 270600 259500 270602
rect 259408 270544 259458 270600
rect 259408 270542 259500 270544
rect 259453 270540 259500 270542
rect 259564 270540 259570 270604
rect 260833 270602 260899 270605
rect 262070 270602 262076 270604
rect 260833 270600 262076 270602
rect 260833 270544 260838 270600
rect 260894 270544 262076 270600
rect 260833 270542 262076 270544
rect 259453 270539 259519 270540
rect 260833 270539 260899 270542
rect 262070 270540 262076 270542
rect 262140 270540 262146 270604
rect 262213 270602 262279 270605
rect 262806 270602 262812 270604
rect 262213 270600 262812 270602
rect 262213 270544 262218 270600
rect 262274 270544 262812 270600
rect 262213 270542 262812 270544
rect 262213 270539 262279 270542
rect 262806 270540 262812 270542
rect 262876 270540 262882 270604
rect 263593 270602 263659 270605
rect 263910 270602 263916 270604
rect 263593 270600 263916 270602
rect 263593 270544 263598 270600
rect 263654 270544 263916 270600
rect 263593 270542 263916 270544
rect 263593 270539 263659 270542
rect 263910 270540 263916 270542
rect 263980 270540 263986 270604
rect 266353 270602 266419 270605
rect 267590 270602 267596 270604
rect 266353 270600 267596 270602
rect 266353 270544 266358 270600
rect 266414 270544 267596 270600
rect 266353 270542 267596 270544
rect 266353 270539 266419 270542
rect 267590 270540 267596 270542
rect 267660 270540 267666 270604
rect 268193 270602 268259 270605
rect 397453 270604 397519 270605
rect 268694 270602 268700 270604
rect 268193 270600 268700 270602
rect 268193 270544 268198 270600
rect 268254 270544 268700 270600
rect 268193 270542 268700 270544
rect 268193 270539 268259 270542
rect 268694 270540 268700 270542
rect 268764 270540 268770 270604
rect 397453 270602 397500 270604
rect 397408 270600 397500 270602
rect 397408 270544 397458 270600
rect 397408 270542 397500 270544
rect 397453 270540 397500 270542
rect 397564 270540 397570 270604
rect 398833 270602 398899 270605
rect 399518 270602 399524 270604
rect 398833 270600 399524 270602
rect 398833 270544 398838 270600
rect 398894 270544 399524 270600
rect 398833 270542 399524 270544
rect 397453 270539 397519 270540
rect 398833 270539 398899 270542
rect 399518 270540 399524 270542
rect 399588 270540 399594 270604
rect 400213 270602 400279 270605
rect 402973 270604 403039 270605
rect 400438 270602 400444 270604
rect 400213 270600 400444 270602
rect 400213 270544 400218 270600
rect 400274 270544 400444 270600
rect 400213 270542 400444 270544
rect 400213 270539 400279 270542
rect 400438 270540 400444 270542
rect 400508 270540 400514 270604
rect 402973 270600 403020 270604
rect 403084 270602 403090 270604
rect 403617 270602 403683 270605
rect 404118 270602 404124 270604
rect 402973 270544 402978 270600
rect 402973 270540 403020 270544
rect 403084 270542 403130 270602
rect 403617 270600 404124 270602
rect 403617 270544 403622 270600
rect 403678 270544 404124 270600
rect 403617 270542 404124 270544
rect 403084 270540 403090 270542
rect 402973 270539 403039 270540
rect 403617 270539 403683 270542
rect 404118 270540 404124 270542
rect 404188 270540 404194 270604
rect 404353 270602 404419 270605
rect 405038 270602 405044 270604
rect 404353 270600 405044 270602
rect 404353 270544 404358 270600
rect 404414 270544 405044 270600
rect 404353 270542 405044 270544
rect 404353 270539 404419 270542
rect 405038 270540 405044 270542
rect 405108 270540 405114 270604
rect 407113 270602 407179 270605
rect 407614 270602 407620 270604
rect 407113 270600 407620 270602
rect 407113 270544 407118 270600
rect 407174 270544 407620 270600
rect 407113 270542 407620 270544
rect 407113 270539 407179 270542
rect 407614 270540 407620 270542
rect 407684 270540 407690 270604
rect 408493 270602 408559 270605
rect 408718 270602 408724 270604
rect 408493 270600 408724 270602
rect 408493 270544 408498 270600
rect 408554 270544 408724 270600
rect 408493 270542 408724 270544
rect 408493 270539 408559 270542
rect 408718 270540 408724 270542
rect 408788 270540 408794 270604
rect 409873 270602 409939 270605
rect 410006 270602 410012 270604
rect 409873 270600 410012 270602
rect 409873 270544 409878 270600
rect 409934 270544 410012 270600
rect 409873 270542 410012 270544
rect 409873 270539 409939 270542
rect 410006 270540 410012 270542
rect 410076 270540 410082 270604
rect 411253 270602 411319 270605
rect 412398 270602 412404 270604
rect 411253 270600 412404 270602
rect 411253 270544 411258 270600
rect 411314 270544 412404 270600
rect 411253 270542 412404 270544
rect 411253 270539 411319 270542
rect 412398 270540 412404 270542
rect 412468 270540 412474 270604
rect 413001 270602 413067 270605
rect 413318 270602 413324 270604
rect 413001 270600 413324 270602
rect 413001 270544 413006 270600
rect 413062 270544 413324 270600
rect 413001 270542 413324 270544
rect 413001 270539 413067 270542
rect 413318 270540 413324 270542
rect 413388 270540 413394 270604
rect 414013 270602 414079 270605
rect 414422 270602 414428 270604
rect 414013 270600 414428 270602
rect 414013 270544 414018 270600
rect 414074 270544 414428 270600
rect 414013 270542 414428 270544
rect 414013 270539 414079 270542
rect 414422 270540 414428 270542
rect 414492 270540 414498 270604
rect 416773 270602 416839 270605
rect 418153 270604 418219 270605
rect 416998 270602 417004 270604
rect 416773 270600 417004 270602
rect 416773 270544 416778 270600
rect 416834 270544 417004 270600
rect 416773 270542 417004 270544
rect 416773 270539 416839 270542
rect 416998 270540 417004 270542
rect 417068 270540 417074 270604
rect 418102 270540 418108 270604
rect 418172 270602 418219 270604
rect 419533 270602 419599 270605
rect 420678 270602 420684 270604
rect 418172 270600 418264 270602
rect 418214 270544 418264 270600
rect 418172 270542 418264 270544
rect 419533 270600 420684 270602
rect 419533 270544 419538 270600
rect 419594 270544 420684 270600
rect 419533 270542 420684 270544
rect 418172 270540 418219 270542
rect 418153 270539 418219 270540
rect 419533 270539 419599 270542
rect 420678 270540 420684 270542
rect 420748 270540 420754 270604
rect 420913 270602 420979 270605
rect 421782 270602 421788 270604
rect 420913 270600 421788 270602
rect 420913 270544 420918 270600
rect 420974 270544 421788 270600
rect 420913 270542 421788 270544
rect 420913 270539 420979 270542
rect 421782 270540 421788 270542
rect 421852 270540 421858 270604
rect 53281 270466 53347 270469
rect 57462 270466 57468 270468
rect 53281 270464 57468 270466
rect 53281 270408 53286 270464
rect 53342 270408 57468 270464
rect 53281 270406 57468 270408
rect 53281 270403 53347 270406
rect 57462 270404 57468 270406
rect 57532 270466 57538 270468
rect 91502 270466 91508 270468
rect 57532 270406 91508 270466
rect 57532 270404 57538 270406
rect 91502 270404 91508 270406
rect 91572 270404 91578 270468
rect 211521 270466 211587 270469
rect 323342 270466 323348 270468
rect 211521 270464 323348 270466
rect 211521 270408 211526 270464
rect 211582 270408 323348 270464
rect 211521 270406 323348 270408
rect 211521 270403 211587 270406
rect 323342 270404 323348 270406
rect 323412 270404 323418 270468
rect 378685 270466 378751 270469
rect 379697 270466 379763 270469
rect 419206 270466 419212 270468
rect 378685 270464 379763 270466
rect 378685 270408 378690 270464
rect 378746 270408 379702 270464
rect 379758 270408 379763 270464
rect 378685 270406 379763 270408
rect 378685 270403 378751 270406
rect 379697 270403 379763 270406
rect 383610 270406 419212 270466
rect 207565 270330 207631 270333
rect 208301 270330 208367 270333
rect 241646 270330 241652 270332
rect 207565 270328 241652 270330
rect 207565 270272 207570 270328
rect 207626 270272 208306 270328
rect 208362 270272 241652 270328
rect 207565 270270 241652 270272
rect 207565 270267 207631 270270
rect 208301 270267 208367 270270
rect 241646 270268 241652 270270
rect 241716 270268 241722 270332
rect 376477 270330 376543 270333
rect 383610 270330 383670 270406
rect 419206 270404 419212 270406
rect 419276 270404 419282 270468
rect 376477 270328 383670 270330
rect 376477 270272 376482 270328
rect 376538 270272 383670 270328
rect 376477 270270 383670 270272
rect 376477 270267 376543 270270
rect 210877 270194 210943 270197
rect 214925 270194 214991 270197
rect 240542 270194 240548 270196
rect 210877 270192 240548 270194
rect 210877 270136 210882 270192
rect 210938 270136 214930 270192
rect 214986 270136 240548 270192
rect 210877 270134 240548 270136
rect 210877 270131 210943 270134
rect 214925 270131 214991 270134
rect 240542 270132 240548 270134
rect 240612 270132 240618 270196
rect 217542 269860 217548 269924
rect 217612 269922 217618 269924
rect 219065 269922 219131 269925
rect 217612 269920 219131 269922
rect 217612 269864 219070 269920
rect 219126 269864 219131 269920
rect 217612 269862 219131 269864
rect 217612 269860 217618 269862
rect 219065 269859 219131 269862
rect 371693 269922 371759 269925
rect 379237 269922 379303 269925
rect 371693 269920 379303 269922
rect 371693 269864 371698 269920
rect 371754 269864 379242 269920
rect 379298 269864 379303 269920
rect 371693 269862 379303 269864
rect 371693 269859 371759 269862
rect 379237 269859 379303 269862
rect 208853 269786 208919 269789
rect 212349 269786 212415 269789
rect 239254 269786 239260 269788
rect 208853 269784 239260 269786
rect 208853 269728 208858 269784
rect 208914 269728 212354 269784
rect 212410 269728 239260 269784
rect 208853 269726 239260 269728
rect 208853 269723 208919 269726
rect 212349 269723 212415 269726
rect 239254 269724 239260 269726
rect 239324 269724 239330 269788
rect 379697 269786 379763 269789
rect 426382 269786 426388 269788
rect 379697 269784 426388 269786
rect 379697 269728 379702 269784
rect 379758 269728 426388 269784
rect 379697 269726 426388 269728
rect 379697 269723 379763 269726
rect 426382 269724 426388 269726
rect 426452 269724 426458 269788
rect 379237 269378 379303 269381
rect 390553 269378 390619 269381
rect 379237 269376 390619 269378
rect 379237 269320 379242 269376
rect 379298 269320 390558 269376
rect 390614 269320 390619 269376
rect 379237 269318 390619 269320
rect 379237 269315 379303 269318
rect 390553 269315 390619 269318
rect 372981 269242 373047 269245
rect 373533 269242 373599 269245
rect 388437 269242 388503 269245
rect 372981 269240 388503 269242
rect 372981 269184 372986 269240
rect 373042 269184 373538 269240
rect 373594 269184 388442 269240
rect 388498 269184 388503 269240
rect 372981 269182 388503 269184
rect 372981 269179 373047 269182
rect 373533 269179 373599 269182
rect 388437 269179 388503 269182
rect 44766 269044 44772 269108
rect 44836 269106 44842 269108
rect 59353 269106 59419 269109
rect 44836 269104 59419 269106
rect 44836 269048 59358 269104
rect 59414 269048 59419 269104
rect 44836 269046 59419 269048
rect 44836 269044 44842 269046
rect 59353 269043 59419 269046
rect 44950 268908 44956 268972
rect 45020 268970 45026 268972
rect 57237 268970 57303 268973
rect 45020 268968 57303 268970
rect 45020 268912 57242 268968
rect 57298 268912 57303 268968
rect 45020 268910 57303 268912
rect 45020 268908 45026 268910
rect 57237 268907 57303 268910
rect 217225 268700 217291 268701
rect 217174 268698 217180 268700
rect 217134 268638 217180 268698
rect 217244 268696 217291 268700
rect 217286 268640 217291 268696
rect 217174 268636 217180 268638
rect 217244 268636 217291 268640
rect 217225 268635 217291 268636
rect -960 267052 480 267292
rect 377990 264964 377996 265028
rect 378060 265026 378066 265028
rect 379053 265026 379119 265029
rect 378060 265024 379119 265026
rect 378060 264968 379058 265024
rect 379114 264968 379119 265024
rect 378060 264966 379119 264968
rect 378060 264964 378066 264966
rect 379053 264963 379119 264966
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect -960 254086 6930 254146
rect -960 253996 480 254086
rect 6870 254010 6930 254086
rect 54334 254010 54340 254012
rect 6870 253950 54340 254010
rect 54334 253948 54340 253950
rect 54404 253948 54410 254012
rect 339718 253404 339724 253468
rect 339788 253466 339794 253468
rect 340781 253466 340847 253469
rect 339788 253464 340847 253466
rect 339788 253408 340786 253464
rect 340842 253408 340847 253464
rect 339788 253406 340847 253408
rect 339788 253404 339794 253406
rect 340781 253403 340847 253406
rect 179638 253268 179644 253332
rect 179708 253330 179714 253332
rect 180149 253330 180215 253333
rect 179708 253328 180215 253330
rect 179708 253272 180154 253328
rect 180210 253272 180215 253328
rect 179708 253270 180215 253272
rect 179708 253268 179714 253270
rect 180149 253267 180215 253270
rect 499798 253268 499804 253332
rect 499868 253330 499874 253332
rect 500861 253330 500927 253333
rect 499868 253328 500927 253330
rect 499868 253272 500866 253328
rect 500922 253272 500927 253328
rect 499868 253270 500927 253272
rect 499868 253268 499874 253270
rect 500861 253267 500927 253270
rect 178534 253132 178540 253196
rect 178604 253194 178610 253196
rect 179321 253194 179387 253197
rect 178604 253192 179387 253194
rect 178604 253136 179326 253192
rect 179382 253136 179387 253192
rect 178604 253134 179387 253136
rect 178604 253132 178610 253134
rect 179321 253131 179387 253134
rect 190862 253132 190868 253196
rect 190932 253194 190938 253196
rect 191741 253194 191807 253197
rect 190932 253192 191807 253194
rect 190932 253136 191746 253192
rect 191802 253136 191807 253192
rect 190932 253134 191807 253136
rect 190932 253132 190938 253134
rect 191741 253131 191807 253134
rect 350942 253132 350948 253196
rect 351012 253194 351018 253196
rect 351821 253194 351887 253197
rect 351012 253192 351887 253194
rect 351012 253136 351826 253192
rect 351882 253136 351887 253192
rect 351012 253134 351887 253136
rect 351012 253132 351018 253134
rect 351821 253131 351887 253134
rect 338430 252996 338436 253060
rect 338500 253058 338506 253060
rect 339401 253058 339467 253061
rect 338500 253056 339467 253058
rect 338500 253000 339406 253056
rect 339462 253000 339467 253056
rect 338500 252998 339467 253000
rect 338500 252996 338506 252998
rect 339401 252995 339467 252998
rect 498510 252724 498516 252788
rect 498580 252786 498586 252788
rect 499205 252786 499271 252789
rect 498580 252784 499271 252786
rect 498580 252728 499210 252784
rect 499266 252728 499271 252784
rect 498580 252726 499271 252728
rect 498580 252724 498586 252726
rect 499205 252723 499271 252726
rect 510889 252652 510955 252653
rect 510838 252650 510844 252652
rect 510798 252590 510844 252650
rect 510908 252648 510955 252652
rect 510950 252592 510955 252648
rect 510838 252588 510844 252590
rect 510908 252588 510955 252592
rect 510889 252587 510955 252588
rect 377397 252514 377463 252517
rect 377990 252514 377996 252516
rect 377397 252512 377996 252514
rect 377397 252456 377402 252512
rect 377458 252456 377996 252512
rect 377397 252454 377996 252456
rect 377397 252451 377463 252454
rect 377990 252452 377996 252454
rect 378060 252452 378066 252516
rect 198825 246258 198891 246261
rect 358905 246258 358971 246261
rect 519077 246258 519143 246261
rect 196558 246256 198891 246258
rect 196558 246200 198830 246256
rect 198886 246200 198891 246256
rect 196558 246198 198891 246200
rect 196558 246190 196618 246198
rect 198825 246195 198891 246198
rect 356562 246256 358971 246258
rect 356562 246200 358910 246256
rect 358966 246200 358971 246256
rect 356562 246198 358971 246200
rect 356562 246190 356622 246198
rect 358905 246195 358971 246198
rect 516558 246256 519143 246258
rect 516558 246200 519082 246256
rect 519138 246200 519143 246256
rect 516558 246198 519143 246200
rect 516558 246190 516618 246198
rect 519077 246195 519143 246198
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect 57145 204234 57211 204237
rect 57513 204234 57579 204237
rect 377029 204234 377095 204237
rect 377305 204234 377371 204237
rect 57145 204232 60062 204234
rect 57145 204176 57150 204232
rect 57206 204176 57518 204232
rect 57574 204176 60062 204232
rect 57145 204174 60062 204176
rect 57145 204171 57211 204174
rect 57513 204171 57579 204174
rect 60002 203894 60062 204174
rect 377029 204232 377371 204234
rect 377029 204176 377034 204232
rect 377090 204176 377310 204232
rect 377366 204176 377371 204232
rect 377029 204174 377371 204176
rect 377029 204171 377095 204174
rect 377305 204171 377371 204174
rect 217409 203962 217475 203965
rect 217593 203962 217659 203965
rect 376937 203962 377003 203965
rect 377305 203962 377371 203965
rect 217409 203960 219450 203962
rect 217409 203904 217414 203960
rect 217470 203904 217598 203960
rect 217654 203924 219450 203960
rect 376937 203960 379530 203962
rect 217654 203904 220064 203924
rect 217409 203902 220064 203904
rect 217409 203899 217475 203902
rect 217593 203899 217659 203902
rect 219390 203864 220064 203902
rect 376937 203904 376942 203960
rect 376998 203904 377310 203960
rect 377366 203924 379530 203960
rect 377366 203904 380052 203924
rect 376937 203902 380052 203904
rect 376937 203899 377003 203902
rect 377305 203899 377371 203902
rect 379470 203864 380052 203902
rect 56777 203554 56843 203557
rect 57329 203554 57395 203557
rect 56777 203552 60062 203554
rect 56777 203496 56782 203552
rect 56838 203496 57334 203552
rect 57390 203496 60062 203552
rect 56777 203494 60062 203496
rect 56777 203491 56843 203494
rect 57329 203491 57395 203494
rect 60002 202942 60062 203494
rect 217133 203010 217199 203013
rect 217593 203010 217659 203013
rect 377029 203010 377095 203013
rect 217133 203008 219450 203010
rect 217133 202952 217138 203008
rect 217194 202952 217598 203008
rect 217654 202972 219450 203008
rect 377029 203008 379530 203010
rect 217654 202952 220064 202972
rect 217133 202950 220064 202952
rect 217133 202947 217199 202950
rect 217593 202947 217659 202950
rect 219390 202912 220064 202950
rect 377029 202952 377034 203008
rect 377090 202972 379530 203008
rect 377090 202952 380052 202972
rect 377029 202950 380052 202952
rect 377029 202947 377095 202950
rect 379470 202912 380052 202950
rect -960 201922 480 202012
rect -960 201862 6930 201922
rect -960 201772 480 201862
rect 6870 201514 6930 201862
rect 53046 201514 53052 201516
rect 6870 201454 53052 201514
rect 53046 201452 53052 201454
rect 53116 201452 53122 201516
rect 56869 201378 56935 201381
rect 57605 201378 57671 201381
rect 376937 201378 377003 201381
rect 377673 201378 377739 201381
rect 56869 201376 60062 201378
rect 56869 201320 56874 201376
rect 56930 201320 57610 201376
rect 57666 201320 60062 201376
rect 56869 201318 60062 201320
rect 56869 201315 56935 201318
rect 57605 201315 57671 201318
rect 60002 200766 60062 201318
rect 376937 201376 377739 201378
rect 376937 201320 376942 201376
rect 376998 201320 377678 201376
rect 377734 201320 377739 201376
rect 376937 201318 377739 201320
rect 376937 201315 377003 201318
rect 377673 201315 377739 201318
rect 217685 200834 217751 200837
rect 377673 200834 377739 200837
rect 217685 200832 219450 200834
rect 217685 200776 217690 200832
rect 217746 200796 219450 200832
rect 377673 200832 379530 200834
rect 217746 200776 220064 200796
rect 217685 200774 220064 200776
rect 217685 200771 217751 200774
rect 219390 200736 220064 200774
rect 377673 200776 377678 200832
rect 377734 200796 379530 200832
rect 377734 200776 380052 200796
rect 377673 200774 380052 200776
rect 377673 200771 377739 200774
rect 379470 200736 380052 200774
rect 57789 199882 57855 199885
rect 217501 199882 217567 199885
rect 377857 199882 377923 199885
rect 57789 199880 60062 199882
rect 57789 199824 57794 199880
rect 57850 199824 60062 199880
rect 57789 199822 60062 199824
rect 57789 199819 57855 199822
rect 60002 199814 60062 199822
rect 217501 199880 219450 199882
rect 217501 199824 217506 199880
rect 217562 199844 219450 199880
rect 377857 199880 379530 199882
rect 217562 199824 220064 199844
rect 217501 199822 220064 199824
rect 217501 199819 217567 199822
rect 219390 199784 220064 199822
rect 377857 199824 377862 199880
rect 377918 199844 379530 199880
rect 377918 199824 380052 199844
rect 377857 199822 380052 199824
rect 377857 199819 377923 199822
rect 379470 199784 380052 199822
rect 57329 198794 57395 198797
rect 57789 198794 57855 198797
rect 57329 198792 57855 198794
rect 57329 198736 57334 198792
rect 57390 198736 57794 198792
rect 57850 198736 57855 198792
rect 57329 198734 57855 198736
rect 57329 198731 57395 198734
rect 57789 198731 57855 198734
rect 217225 198794 217291 198797
rect 217501 198794 217567 198797
rect 217225 198792 217567 198794
rect 217225 198736 217230 198792
rect 217286 198736 217506 198792
rect 217562 198736 217567 198792
rect 217225 198734 217567 198736
rect 217225 198731 217291 198734
rect 217501 198731 217567 198734
rect 377213 198794 377279 198797
rect 377857 198794 377923 198797
rect 377213 198792 377923 198794
rect 377213 198736 377218 198792
rect 377274 198736 377862 198792
rect 377918 198736 377923 198792
rect 377213 198734 377923 198736
rect 377213 198731 377279 198734
rect 377857 198731 377923 198734
rect 57789 198114 57855 198117
rect 216765 198114 216831 198117
rect 217501 198114 217567 198117
rect 377673 198114 377739 198117
rect 57789 198112 60062 198114
rect 57789 198056 57794 198112
rect 57850 198056 60062 198112
rect 57789 198054 60062 198056
rect 57789 198051 57855 198054
rect 60002 198046 60062 198054
rect 216765 198112 219450 198114
rect 216765 198056 216770 198112
rect 216826 198056 217506 198112
rect 217562 198076 219450 198112
rect 377673 198112 379530 198114
rect 217562 198056 220064 198076
rect 216765 198054 220064 198056
rect 216765 198051 216831 198054
rect 217501 198051 217567 198054
rect 219390 198016 220064 198054
rect 377673 198056 377678 198112
rect 377734 198076 379530 198112
rect 377734 198056 380052 198076
rect 377673 198054 380052 198056
rect 377673 198051 377739 198054
rect 379470 198016 380052 198054
rect 216765 197026 216831 197029
rect 217777 197026 217843 197029
rect 377581 197026 377647 197029
rect 377857 197026 377923 197029
rect 216765 197024 219450 197026
rect 216765 196968 216770 197024
rect 216826 196968 217782 197024
rect 217838 196988 219450 197024
rect 377581 197024 379530 197026
rect 217838 196968 220064 196988
rect 216765 196966 220064 196968
rect 216765 196963 216831 196966
rect 217777 196963 217843 196966
rect 57421 196346 57487 196349
rect 60002 196346 60062 196958
rect 219390 196928 220064 196966
rect 377581 196968 377586 197024
rect 377642 196968 377862 197024
rect 377918 196988 379530 197024
rect 377918 196968 380052 196988
rect 377581 196966 380052 196968
rect 377581 196963 377647 196966
rect 377857 196963 377923 196966
rect 379470 196928 380052 196966
rect 57421 196344 60062 196346
rect 57421 196288 57426 196344
rect 57482 196288 60062 196344
rect 57421 196286 60062 196288
rect 57421 196283 57487 196286
rect 57053 195258 57119 195261
rect 57697 195258 57763 195261
rect 216949 195258 217015 195261
rect 217777 195258 217843 195261
rect 377121 195258 377187 195261
rect 377765 195258 377831 195261
rect 57053 195256 60062 195258
rect 57053 195200 57058 195256
rect 57114 195200 57702 195256
rect 57758 195200 60062 195256
rect 57053 195198 60062 195200
rect 57053 195195 57119 195198
rect 57697 195195 57763 195198
rect 60002 195190 60062 195198
rect 216949 195256 219450 195258
rect 216949 195200 216954 195256
rect 217010 195200 217782 195256
rect 217838 195220 219450 195256
rect 377121 195256 379530 195258
rect 217838 195200 220064 195220
rect 216949 195198 220064 195200
rect 216949 195195 217015 195198
rect 217777 195195 217843 195198
rect 219390 195160 220064 195198
rect 377121 195200 377126 195256
rect 377182 195200 377770 195256
rect 377826 195220 379530 195256
rect 377826 195200 380052 195220
rect 377121 195198 380052 195200
rect 377121 195195 377187 195198
rect 377765 195195 377831 195198
rect 379470 195160 380052 195198
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 199285 186418 199351 186421
rect 359273 186418 359339 186421
rect 359457 186418 359523 186421
rect 518893 186418 518959 186421
rect 519353 186418 519419 186421
rect 196558 186416 199351 186418
rect 196558 186360 199290 186416
rect 199346 186360 199351 186416
rect 196558 186358 199351 186360
rect 196558 186350 196618 186358
rect 199285 186355 199351 186358
rect 356562 186416 359523 186418
rect 356562 186360 359278 186416
rect 359334 186360 359462 186416
rect 359518 186360 359523 186416
rect 356562 186358 359523 186360
rect 356562 186350 356622 186358
rect 359273 186355 359339 186358
rect 359457 186355 359523 186358
rect 516558 186416 519419 186418
rect 516558 186360 518898 186416
rect 518954 186360 519358 186416
rect 519414 186360 519419 186416
rect 516558 186358 519419 186360
rect 516558 186350 516618 186358
rect 518893 186355 518959 186358
rect 519353 186355 519419 186358
rect 198917 184922 198983 184925
rect 199193 184922 199259 184925
rect 358813 184922 358879 184925
rect 359365 184922 359431 184925
rect 196558 184920 199259 184922
rect 196558 184864 198922 184920
rect 198978 184864 199198 184920
rect 199254 184864 199259 184920
rect 196558 184862 199259 184864
rect 196558 184718 196618 184862
rect 198917 184859 198983 184862
rect 199193 184859 199259 184862
rect 356562 184920 359431 184922
rect 356562 184864 358818 184920
rect 358874 184864 359370 184920
rect 359426 184864 359431 184920
rect 356562 184862 359431 184864
rect 356562 184718 356622 184862
rect 358813 184859 358879 184862
rect 359365 184859 359431 184862
rect 519445 184786 519511 184789
rect 520181 184786 520247 184789
rect 516558 184784 520247 184786
rect 516558 184728 519450 184784
rect 519506 184728 520186 184784
rect 520242 184728 520247 184784
rect 516558 184726 520247 184728
rect 516558 184718 516618 184726
rect 519445 184723 519511 184726
rect 520181 184723 520247 184726
rect 198733 183562 198799 183565
rect 198917 183562 198983 183565
rect 196558 183560 198983 183562
rect 196558 183504 198738 183560
rect 198794 183504 198922 183560
rect 198978 183504 198983 183560
rect 196558 183502 198983 183504
rect 196558 183358 196618 183502
rect 198733 183499 198799 183502
rect 198917 183499 198983 183502
rect 359181 183426 359247 183429
rect 518985 183426 519051 183429
rect 519353 183426 519419 183429
rect 520089 183426 520155 183429
rect 356562 183424 359247 183426
rect 356562 183368 359186 183424
rect 359242 183368 359247 183424
rect 356562 183366 359247 183368
rect 356562 183358 356622 183366
rect 359181 183363 359247 183366
rect 516558 183424 520155 183426
rect 516558 183368 518990 183424
rect 519046 183368 519358 183424
rect 519414 183368 520094 183424
rect 520150 183368 520155 183424
rect 516558 183366 520155 183368
rect 516558 183358 516618 183366
rect 518985 183363 519051 183366
rect 519353 183363 519419 183366
rect 520089 183363 520155 183366
rect 198733 182066 198799 182069
rect 199009 182066 199075 182069
rect 359089 182066 359155 182069
rect 359549 182066 359615 182069
rect 196558 182064 199075 182066
rect 196558 182008 198738 182064
rect 198794 182008 199014 182064
rect 199070 182008 199075 182064
rect 196558 182006 199075 182008
rect 196558 181862 196618 182006
rect 198733 182003 198799 182006
rect 199009 182003 199075 182006
rect 356562 182064 359615 182066
rect 356562 182008 359094 182064
rect 359150 182008 359554 182064
rect 359610 182008 359615 182064
rect 356562 182006 359615 182008
rect 356562 181862 356622 182006
rect 359089 182003 359155 182006
rect 359549 182003 359615 182006
rect 518985 181930 519051 181933
rect 519169 181930 519235 181933
rect 516558 181928 519235 181930
rect 516558 181872 518990 181928
rect 519046 181872 519174 181928
rect 519230 181872 519235 181928
rect 516558 181870 519235 181872
rect 516558 181862 516618 181870
rect 518985 181867 519051 181870
rect 519169 181867 519235 181870
rect 199101 180706 199167 180709
rect 358997 180706 359063 180709
rect 519261 180706 519327 180709
rect 196558 180704 199167 180706
rect 196558 180648 199106 180704
rect 199162 180648 199167 180704
rect 196558 180646 199167 180648
rect 196558 180638 196618 180646
rect 199101 180643 199167 180646
rect 356562 180704 359063 180706
rect 356562 180648 359002 180704
rect 359058 180648 359063 180704
rect 356562 180646 359063 180648
rect 356562 180638 356622 180646
rect 358997 180643 359063 180646
rect 516558 180704 519327 180706
rect 516558 180648 519266 180704
rect 519322 180648 519327 180704
rect 516558 180646 519327 180648
rect 516558 180638 516618 180646
rect 519261 180643 519327 180646
rect 358997 179482 359063 179485
rect 359273 179482 359339 179485
rect 358997 179480 359339 179482
rect 358997 179424 359002 179480
rect 359058 179424 359278 179480
rect 359334 179424 359339 179480
rect 358997 179422 359339 179424
rect 358997 179419 359063 179422
rect 359273 179419 359339 179422
rect 583520 179060 584960 179300
rect 58893 177578 58959 177581
rect 58893 177576 60062 177578
rect 58893 177520 58898 177576
rect 58954 177520 60062 177576
rect 58893 177518 60062 177520
rect 58893 177515 58959 177518
rect 60002 176966 60062 177518
rect 216673 177034 216739 177037
rect 376937 177034 377003 177037
rect 216673 177032 219450 177034
rect 216673 176976 216678 177032
rect 216734 176996 219450 177032
rect 376937 177032 379530 177034
rect 216734 176976 220064 176996
rect 216673 176974 220064 176976
rect 216673 176971 216739 176974
rect 219390 176936 220064 176974
rect 376937 176976 376942 177032
rect 376998 176996 379530 177032
rect 376998 176976 380052 176996
rect 376937 176974 380052 176976
rect 376937 176971 377003 176974
rect 379470 176936 380052 176974
rect -960 175796 480 176036
rect 57462 175884 57468 175948
rect 57532 175946 57538 175948
rect 59445 175946 59511 175949
rect 57532 175944 59511 175946
rect 57532 175888 59450 175944
rect 59506 175888 59511 175944
rect 57532 175886 59511 175888
rect 57532 175884 57538 175886
rect 59445 175883 59511 175886
rect 57881 175810 57947 175813
rect 57881 175808 60062 175810
rect 57881 175752 57886 175808
rect 57942 175752 60062 175808
rect 57881 175750 60062 175752
rect 57881 175747 57947 175750
rect 60002 175334 60062 175750
rect 216673 175402 216739 175405
rect 376937 175402 377003 175405
rect 216673 175400 219450 175402
rect 216673 175344 216678 175400
rect 216734 175364 219450 175400
rect 376937 175400 379530 175402
rect 216734 175344 220064 175364
rect 216673 175342 220064 175344
rect 216673 175339 216739 175342
rect 219390 175304 220064 175342
rect 376937 175344 376942 175400
rect 376998 175364 379530 175400
rect 376998 175344 380052 175364
rect 376937 175342 380052 175344
rect 376937 175339 377003 175342
rect 379470 175304 380052 175342
rect 57646 175068 57652 175132
rect 57716 175130 57722 175132
rect 216949 175130 217015 175133
rect 376937 175130 377003 175133
rect 57716 175092 59554 175130
rect 216949 175128 219450 175130
rect 57716 175070 60032 175092
rect 57716 175068 57722 175070
rect 59494 175032 60032 175070
rect 216949 175072 216954 175128
rect 217010 175092 219450 175128
rect 376937 175128 379530 175130
rect 217010 175072 220064 175092
rect 216949 175070 220064 175072
rect 216949 175067 217015 175070
rect 219390 175032 220064 175070
rect 376937 175072 376942 175128
rect 376998 175092 379530 175128
rect 376998 175072 380052 175092
rect 376937 175070 380052 175072
rect 376937 175067 377003 175070
rect 379470 175032 380052 175070
rect 57830 166908 57836 166972
rect 57900 166970 57906 166972
rect 57900 166910 143572 166970
rect 57900 166908 57906 166910
rect 96061 166836 96127 166837
rect 98453 166836 98519 166837
rect 101029 166836 101095 166837
rect 105813 166836 105879 166837
rect 108205 166836 108271 166837
rect 138473 166836 138539 166837
rect 140865 166836 140931 166837
rect 143512 166836 143572 166910
rect 202270 166908 202276 166972
rect 202340 166970 202346 166972
rect 202340 166910 313500 166970
rect 202340 166908 202346 166910
rect 145925 166836 145991 166837
rect 313440 166836 313500 166910
rect 356646 166908 356652 166972
rect 356716 166970 356722 166972
rect 356716 166910 471052 166970
rect 356716 166908 356722 166910
rect 418429 166836 418495 166837
rect 421005 166836 421071 166837
rect 428273 166836 428339 166837
rect 430941 166836 431007 166837
rect 433609 166836 433675 166837
rect 470992 166836 471052 166910
rect 473445 166836 473511 166837
rect 47894 166772 47900 166836
rect 47964 166834 47970 166836
rect 93710 166834 93716 166836
rect 47964 166774 93716 166834
rect 47964 166772 47970 166774
rect 93710 166772 93716 166774
rect 93780 166772 93786 166836
rect 96061 166834 96108 166836
rect 96016 166832 96108 166834
rect 96016 166776 96066 166832
rect 96016 166774 96108 166776
rect 96061 166772 96108 166774
rect 96172 166772 96178 166836
rect 98453 166834 98500 166836
rect 98408 166832 98500 166834
rect 98408 166776 98458 166832
rect 98408 166774 98500 166776
rect 98453 166772 98500 166774
rect 98564 166772 98570 166836
rect 101029 166834 101076 166836
rect 100984 166832 101076 166834
rect 100984 166776 101034 166832
rect 100984 166774 101076 166776
rect 101029 166772 101076 166774
rect 101140 166772 101146 166836
rect 105813 166834 105860 166836
rect 105768 166832 105860 166834
rect 105768 166776 105818 166832
rect 105768 166774 105860 166776
rect 105813 166772 105860 166774
rect 105924 166772 105930 166836
rect 108205 166834 108252 166836
rect 108160 166832 108252 166834
rect 108160 166776 108210 166832
rect 108160 166774 108252 166776
rect 108205 166772 108252 166774
rect 108316 166772 108322 166836
rect 138472 166772 138478 166836
rect 138542 166834 138548 166836
rect 138542 166774 138630 166834
rect 140865 166832 140926 166836
rect 140865 166776 140870 166832
rect 138542 166772 138548 166774
rect 140865 166772 140926 166776
rect 140990 166834 140996 166836
rect 140990 166774 141022 166834
rect 140990 166772 140996 166774
rect 143504 166772 143510 166836
rect 143574 166772 143580 166836
rect 145925 166832 145958 166836
rect 146022 166834 146028 166836
rect 145925 166776 145930 166832
rect 145925 166772 145958 166776
rect 146022 166774 146082 166834
rect 146022 166772 146028 166774
rect 202454 166772 202460 166836
rect 202524 166834 202530 166836
rect 305952 166834 305958 166836
rect 202524 166774 305958 166834
rect 202524 166772 202530 166774
rect 305952 166772 305958 166774
rect 306022 166772 306028 166836
rect 313432 166772 313438 166836
rect 313502 166772 313508 166836
rect 418429 166834 418476 166836
rect 418384 166832 418476 166834
rect 418384 166776 418434 166832
rect 418384 166774 418476 166776
rect 418429 166772 418476 166774
rect 418540 166772 418546 166836
rect 421005 166834 421052 166836
rect 420960 166832 421052 166834
rect 420960 166776 421010 166832
rect 420960 166774 421052 166776
rect 421005 166772 421052 166774
rect 421116 166772 421122 166836
rect 428273 166832 428286 166836
rect 428350 166834 428356 166836
rect 428273 166776 428278 166832
rect 428273 166772 428286 166776
rect 428350 166774 428430 166834
rect 430941 166832 431006 166836
rect 430941 166776 430946 166832
rect 431002 166776 431006 166832
rect 428350 166772 428356 166774
rect 430941 166772 431006 166776
rect 431070 166834 431076 166836
rect 433584 166834 433590 166836
rect 431070 166774 431098 166834
rect 433518 166774 433590 166834
rect 433654 166832 433675 166836
rect 433670 166776 433675 166832
rect 431070 166772 431076 166774
rect 433584 166772 433590 166774
rect 433654 166772 433675 166776
rect 470984 166772 470990 166836
rect 471054 166772 471060 166836
rect 473432 166834 473438 166836
rect 473354 166774 473438 166834
rect 473502 166832 473511 166836
rect 473506 166776 473511 166832
rect 473432 166772 473438 166774
rect 473502 166772 473511 166776
rect 96061 166771 96127 166772
rect 98453 166771 98519 166772
rect 101029 166771 101095 166772
rect 105813 166771 105879 166772
rect 108205 166771 108271 166772
rect 138473 166771 138539 166772
rect 140865 166771 140931 166772
rect 145925 166771 145991 166772
rect 418429 166771 418495 166772
rect 421005 166771 421071 166772
rect 428273 166771 428339 166772
rect 430941 166771 431007 166772
rect 433609 166771 433675 166772
rect 473445 166771 473511 166772
rect 475837 166836 475903 166837
rect 478413 166836 478479 166837
rect 480897 166836 480963 166837
rect 475837 166832 475886 166836
rect 475950 166834 475956 166836
rect 475837 166776 475842 166832
rect 475837 166772 475886 166776
rect 475950 166774 475994 166834
rect 478413 166832 478470 166836
rect 478534 166834 478540 166836
rect 478413 166776 478418 166832
rect 475950 166772 475956 166774
rect 478413 166772 478470 166776
rect 478534 166774 478570 166834
rect 480897 166832 480918 166836
rect 480982 166834 480988 166836
rect 480897 166776 480902 166832
rect 478534 166772 478540 166774
rect 480897 166772 480918 166776
rect 480982 166774 481054 166834
rect 480982 166772 480988 166774
rect 475837 166771 475903 166772
rect 478413 166771 478479 166772
rect 480897 166771 480963 166772
rect 163313 166700 163379 166701
rect 163313 166696 163366 166700
rect 163430 166698 163436 166700
rect 163313 166640 163318 166696
rect 163313 166636 163366 166640
rect 163430 166638 163470 166698
rect 163430 166636 163436 166638
rect 203006 166636 203012 166700
rect 203076 166698 203082 166700
rect 288065 166698 288131 166701
rect 203076 166696 288131 166698
rect 203076 166640 288070 166696
rect 288126 166640 288131 166696
rect 203076 166638 288131 166640
rect 203076 166636 203082 166638
rect 163313 166635 163379 166636
rect 288065 166635 288131 166638
rect 288249 166700 288315 166701
rect 291009 166700 291075 166701
rect 483381 166700 483447 166701
rect 485957 166700 486023 166701
rect 288249 166696 288278 166700
rect 288342 166698 288348 166700
rect 290992 166698 290998 166700
rect 288249 166640 288254 166696
rect 288249 166636 288278 166640
rect 288342 166638 288406 166698
rect 290918 166638 290998 166698
rect 291062 166696 291075 166700
rect 483360 166698 483366 166700
rect 291070 166640 291075 166696
rect 288342 166636 288348 166638
rect 290992 166636 290998 166638
rect 291062 166636 291075 166640
rect 483290 166638 483366 166698
rect 483430 166696 483447 166700
rect 485944 166698 485950 166700
rect 483442 166640 483447 166696
rect 483360 166636 483366 166638
rect 483430 166636 483447 166640
rect 485866 166638 485950 166698
rect 486014 166696 486023 166700
rect 486018 166640 486023 166696
rect 485944 166636 485950 166638
rect 486014 166636 486023 166640
rect 288249 166635 288315 166636
rect 291009 166635 291075 166636
rect 483381 166635 483447 166636
rect 485957 166635 486023 166636
rect 111149 166564 111215 166565
rect 111136 166562 111142 166564
rect 111058 166502 111142 166562
rect 111206 166560 111215 166564
rect 111210 166504 111215 166560
rect 111136 166500 111142 166502
rect 111206 166500 111215 166504
rect 111149 166499 111215 166500
rect 116945 166564 117011 166565
rect 148501 166564 148567 166565
rect 434345 166564 434411 166565
rect 503253 166564 503319 166565
rect 116945 166560 116990 166564
rect 117054 166562 117060 166564
rect 148501 166562 148548 166564
rect 116945 166504 116950 166560
rect 116945 166500 116990 166504
rect 117054 166502 117102 166562
rect 148456 166560 148548 166562
rect 148456 166504 148506 166560
rect 148456 166502 148548 166504
rect 117054 166500 117060 166502
rect 148501 166500 148548 166502
rect 148612 166500 148618 166564
rect 213494 166500 213500 166564
rect 213564 166562 213570 166564
rect 303504 166562 303510 166564
rect 213564 166502 303510 166562
rect 213564 166500 213570 166502
rect 303504 166500 303510 166502
rect 303574 166500 303580 166564
rect 434345 166560 434406 166564
rect 434345 166504 434350 166560
rect 434345 166500 434406 166504
rect 434470 166562 434476 166564
rect 503216 166562 503222 166564
rect 434470 166502 434502 166562
rect 503162 166502 503222 166562
rect 503286 166560 503319 166564
rect 503314 166504 503319 166560
rect 434470 166500 434476 166502
rect 503216 166500 503222 166502
rect 503286 166500 503319 166504
rect 116945 166499 117011 166500
rect 148501 166499 148567 166500
rect 434345 166499 434411 166500
rect 503253 166499 503319 166500
rect 153285 166428 153351 166429
rect 260925 166428 260991 166429
rect 265893 166428 265959 166429
rect 153285 166426 153332 166428
rect 153240 166424 153332 166426
rect 153240 166368 153290 166424
rect 153240 166366 153332 166368
rect 153285 166364 153332 166366
rect 153396 166364 153402 166428
rect 196566 166364 196572 166428
rect 196636 166426 196642 166428
rect 260925 166426 260972 166428
rect 196636 166366 253950 166426
rect 260880 166424 260972 166426
rect 260880 166368 260930 166424
rect 260880 166366 260972 166368
rect 196636 166364 196642 166366
rect 153285 166363 153351 166364
rect 253890 166290 253950 166366
rect 260925 166364 260972 166366
rect 261036 166364 261042 166428
rect 265893 166426 265940 166428
rect 265848 166424 265940 166426
rect 265848 166368 265898 166424
rect 265848 166366 265940 166368
rect 265893 166364 265940 166366
rect 266004 166364 266010 166428
rect 288065 166426 288131 166429
rect 293309 166428 293375 166429
rect 298461 166428 298527 166429
rect 293309 166426 293356 166428
rect 288065 166424 292590 166426
rect 288065 166368 288070 166424
rect 288126 166368 292590 166424
rect 288065 166366 292590 166368
rect 293264 166424 293356 166426
rect 293264 166368 293314 166424
rect 293264 166366 293356 166368
rect 260925 166363 260991 166364
rect 265893 166363 265959 166364
rect 288065 166363 288131 166366
rect 285949 166292 286015 166293
rect 270902 166290 270908 166292
rect 253890 166230 270908 166290
rect 270902 166228 270908 166230
rect 270972 166228 270978 166292
rect 285949 166288 285996 166292
rect 286060 166290 286066 166292
rect 292530 166290 292590 166366
rect 293309 166364 293356 166366
rect 293420 166364 293426 166428
rect 298461 166426 298508 166428
rect 298416 166424 298508 166426
rect 298416 166368 298466 166424
rect 298416 166366 298508 166368
rect 298461 166364 298508 166366
rect 298572 166364 298578 166428
rect 293309 166363 293375 166364
rect 298461 166363 298527 166364
rect 423397 166292 423463 166293
rect 295926 166290 295932 166292
rect 285949 166232 285954 166288
rect 285949 166228 285996 166232
rect 286060 166230 286106 166290
rect 292530 166230 295932 166290
rect 286060 166228 286066 166230
rect 295926 166228 295932 166230
rect 295996 166228 296002 166292
rect 423397 166290 423444 166292
rect 423352 166288 423444 166290
rect 423352 166232 423402 166288
rect 423352 166230 423444 166232
rect 423397 166228 423444 166230
rect 423508 166228 423514 166292
rect 285949 166227 286015 166228
rect 423397 166227 423463 166228
rect 583520 165732 584960 165972
rect 81433 165610 81499 165613
rect 81750 165610 81756 165612
rect 81433 165608 81756 165610
rect 81433 165552 81438 165608
rect 81494 165552 81756 165608
rect 81433 165550 81756 165552
rect 81433 165547 81499 165550
rect 81750 165548 81756 165550
rect 81820 165548 81826 165612
rect 84193 165610 84259 165613
rect 85430 165610 85436 165612
rect 84193 165608 85436 165610
rect 84193 165552 84198 165608
rect 84254 165552 85436 165608
rect 84193 165550 85436 165552
rect 84193 165547 84259 165550
rect 85430 165548 85436 165550
rect 85500 165548 85506 165612
rect 91185 165610 91251 165613
rect 92422 165610 92428 165612
rect 91185 165608 92428 165610
rect 91185 165552 91190 165608
rect 91246 165552 92428 165608
rect 91185 165550 92428 165552
rect 91185 165547 91251 165550
rect 92422 165548 92428 165550
rect 92492 165548 92498 165612
rect 95233 165610 95299 165613
rect 99373 165612 99439 165613
rect 103513 165612 103579 165613
rect 95734 165610 95740 165612
rect 95233 165608 95740 165610
rect 95233 165552 95238 165608
rect 95294 165552 95740 165608
rect 95233 165550 95740 165552
rect 95233 165547 95299 165550
rect 95734 165548 95740 165550
rect 95804 165548 95810 165612
rect 99373 165608 99420 165612
rect 99484 165610 99490 165612
rect 99373 165552 99378 165608
rect 99373 165548 99420 165552
rect 99484 165550 99530 165610
rect 99484 165548 99490 165550
rect 103462 165548 103468 165612
rect 103532 165610 103579 165612
rect 109309 165610 109375 165613
rect 110965 165612 111031 165613
rect 113541 165612 113607 165613
rect 115933 165612 115999 165613
rect 109718 165610 109724 165612
rect 103532 165608 103624 165610
rect 103574 165552 103624 165608
rect 103532 165550 103624 165552
rect 109309 165608 109724 165610
rect 109309 165552 109314 165608
rect 109370 165552 109724 165608
rect 109309 165550 109724 165552
rect 103532 165548 103579 165550
rect 99373 165547 99439 165548
rect 103513 165547 103579 165548
rect 109309 165547 109375 165550
rect 109718 165548 109724 165550
rect 109788 165548 109794 165612
rect 110965 165608 111012 165612
rect 111076 165610 111082 165612
rect 110965 165552 110970 165608
rect 110965 165548 111012 165552
rect 111076 165550 111122 165610
rect 113541 165608 113588 165612
rect 113652 165610 113658 165612
rect 113541 165552 113546 165608
rect 111076 165548 111082 165550
rect 113541 165548 113588 165552
rect 113652 165550 113698 165610
rect 115933 165608 115980 165612
rect 116044 165610 116050 165612
rect 117865 165610 117931 165613
rect 117998 165610 118004 165612
rect 115933 165552 115938 165608
rect 113652 165548 113658 165550
rect 115933 165548 115980 165552
rect 116044 165550 116090 165610
rect 117865 165608 118004 165610
rect 117865 165552 117870 165608
rect 117926 165552 118004 165608
rect 117865 165550 118004 165552
rect 116044 165548 116050 165550
rect 110965 165547 111031 165548
rect 113541 165547 113607 165548
rect 115933 165547 115999 165548
rect 117865 165547 117931 165550
rect 117998 165548 118004 165550
rect 118068 165548 118074 165612
rect 118141 165610 118207 165613
rect 120901 165612 120967 165613
rect 123477 165612 123543 165613
rect 125869 165612 125935 165613
rect 118366 165610 118372 165612
rect 118141 165608 118372 165610
rect 118141 165552 118146 165608
rect 118202 165552 118372 165608
rect 118141 165550 118372 165552
rect 118141 165547 118207 165550
rect 118366 165548 118372 165550
rect 118436 165548 118442 165612
rect 120901 165608 120948 165612
rect 121012 165610 121018 165612
rect 120901 165552 120906 165608
rect 120901 165548 120948 165552
rect 121012 165550 121058 165610
rect 123477 165608 123524 165612
rect 123588 165610 123594 165612
rect 123477 165552 123482 165608
rect 121012 165548 121018 165550
rect 123477 165548 123524 165552
rect 123588 165550 123634 165610
rect 125869 165608 125916 165612
rect 125980 165610 125986 165612
rect 128353 165610 128419 165613
rect 128486 165610 128492 165612
rect 125869 165552 125874 165608
rect 123588 165548 123594 165550
rect 125869 165548 125916 165552
rect 125980 165550 126026 165610
rect 128353 165608 128492 165610
rect 128353 165552 128358 165608
rect 128414 165552 128492 165608
rect 128353 165550 128492 165552
rect 125980 165548 125986 165550
rect 120901 165547 120967 165548
rect 123477 165547 123543 165548
rect 125869 165547 125935 165548
rect 128353 165547 128419 165550
rect 128486 165548 128492 165550
rect 128556 165548 128562 165612
rect 129733 165610 129799 165613
rect 130878 165610 130884 165612
rect 129733 165608 130884 165610
rect 129733 165552 129738 165608
rect 129794 165552 130884 165608
rect 129733 165550 130884 165552
rect 129733 165547 129799 165550
rect 130878 165548 130884 165550
rect 130948 165548 130954 165612
rect 132493 165610 132559 165613
rect 133454 165610 133460 165612
rect 132493 165608 133460 165610
rect 132493 165552 132498 165608
rect 132554 165552 133460 165608
rect 132493 165550 133460 165552
rect 132493 165547 132559 165550
rect 133454 165548 133460 165550
rect 133524 165548 133530 165612
rect 135253 165610 135319 165613
rect 135846 165610 135852 165612
rect 135253 165608 135852 165610
rect 135253 165552 135258 165608
rect 135314 165552 135852 165608
rect 135253 165550 135852 165552
rect 135253 165547 135319 165550
rect 135846 165548 135852 165550
rect 135916 165548 135922 165612
rect 150433 165610 150499 165613
rect 183185 165612 183251 165613
rect 150934 165610 150940 165612
rect 150433 165608 150940 165610
rect 150433 165552 150438 165608
rect 150494 165552 150940 165608
rect 150433 165550 150940 165552
rect 150433 165547 150499 165550
rect 150934 165548 150940 165550
rect 151004 165548 151010 165612
rect 183134 165610 183140 165612
rect 183094 165550 183140 165610
rect 183204 165608 183251 165612
rect 183246 165552 183251 165608
rect 183134 165548 183140 165550
rect 183204 165548 183251 165552
rect 183185 165547 183251 165548
rect 183461 165612 183527 165613
rect 183461 165608 183508 165612
rect 183572 165610 183578 165612
rect 218237 165610 218303 165613
rect 236085 165612 236151 165613
rect 218646 165610 218652 165612
rect 183461 165552 183466 165608
rect 183461 165548 183508 165552
rect 183572 165550 183618 165610
rect 218237 165608 218652 165610
rect 218237 165552 218242 165608
rect 218298 165552 218652 165608
rect 218237 165550 218652 165552
rect 183572 165548 183578 165550
rect 183461 165547 183527 165548
rect 218237 165547 218303 165550
rect 218646 165548 218652 165550
rect 218716 165548 218722 165612
rect 236085 165610 236132 165612
rect 236040 165608 236132 165610
rect 236040 165552 236090 165608
rect 236040 165550 236132 165552
rect 236085 165548 236132 165550
rect 236196 165548 236202 165612
rect 238753 165610 238819 165613
rect 239622 165610 239628 165612
rect 238753 165608 239628 165610
rect 238753 165552 238758 165608
rect 238814 165552 239628 165608
rect 238753 165550 239628 165552
rect 236085 165547 236151 165548
rect 238753 165547 238819 165550
rect 239622 165548 239628 165550
rect 239692 165548 239698 165612
rect 242893 165610 242959 165613
rect 243118 165610 243124 165612
rect 242893 165608 243124 165610
rect 242893 165552 242898 165608
rect 242954 165552 243124 165608
rect 242893 165550 243124 165552
rect 242893 165547 242959 165550
rect 243118 165548 243124 165550
rect 243188 165548 243194 165612
rect 247125 165610 247191 165613
rect 247534 165610 247540 165612
rect 247125 165608 247540 165610
rect 247125 165552 247130 165608
rect 247186 165552 247540 165608
rect 247125 165550 247540 165552
rect 247125 165547 247191 165550
rect 247534 165548 247540 165550
rect 247604 165548 247610 165612
rect 255313 165610 255379 165613
rect 256182 165610 256188 165612
rect 255313 165608 256188 165610
rect 255313 165552 255318 165608
rect 255374 165552 256188 165608
rect 255313 165550 256188 165552
rect 255313 165547 255379 165550
rect 256182 165548 256188 165550
rect 256252 165548 256258 165612
rect 258022 165548 258028 165612
rect 258092 165610 258098 165612
rect 258165 165610 258231 165613
rect 258092 165608 258231 165610
rect 258092 165552 258170 165608
rect 258226 165552 258231 165608
rect 258092 165550 258231 165552
rect 258092 165548 258098 165550
rect 258165 165547 258231 165550
rect 260833 165610 260899 165613
rect 261702 165610 261708 165612
rect 260833 165608 261708 165610
rect 260833 165552 260838 165608
rect 260894 165552 261708 165608
rect 260833 165550 261708 165552
rect 260833 165547 260899 165550
rect 261702 165548 261708 165550
rect 261772 165548 261778 165612
rect 277393 165610 277459 165613
rect 278446 165610 278452 165612
rect 277393 165608 278452 165610
rect 277393 165552 277398 165608
rect 277454 165552 278452 165608
rect 277393 165550 278452 165552
rect 277393 165547 277459 165550
rect 278446 165548 278452 165550
rect 278516 165548 278522 165612
rect 280153 165610 280219 165613
rect 283373 165612 283439 165613
rect 300853 165612 300919 165613
rect 280838 165610 280844 165612
rect 280153 165608 280844 165610
rect 280153 165552 280158 165608
rect 280214 165552 280844 165608
rect 280153 165550 280844 165552
rect 280153 165547 280219 165550
rect 280838 165548 280844 165550
rect 280908 165548 280914 165612
rect 283373 165608 283420 165612
rect 283484 165610 283490 165612
rect 300853 165610 300900 165612
rect 283373 165552 283378 165608
rect 283373 165548 283420 165552
rect 283484 165550 283530 165610
rect 300808 165608 300900 165610
rect 300808 165552 300858 165608
rect 300808 165550 300900 165552
rect 283484 165548 283490 165550
rect 300853 165548 300900 165550
rect 300964 165548 300970 165612
rect 308213 165610 308279 165613
rect 320909 165612 320975 165613
rect 325877 165612 325943 165613
rect 343265 165612 343331 165613
rect 343449 165612 343515 165613
rect 308438 165610 308444 165612
rect 308213 165608 308444 165610
rect 308213 165552 308218 165608
rect 308274 165552 308444 165608
rect 308213 165550 308444 165552
rect 283373 165547 283439 165548
rect 300853 165547 300919 165548
rect 308213 165547 308279 165550
rect 308438 165548 308444 165550
rect 308508 165548 308514 165612
rect 320909 165608 320956 165612
rect 321020 165610 321026 165612
rect 320909 165552 320914 165608
rect 320909 165548 320956 165552
rect 321020 165550 321066 165610
rect 325877 165608 325924 165612
rect 325988 165610 325994 165612
rect 343214 165610 343220 165612
rect 325877 165552 325882 165608
rect 321020 165548 321026 165550
rect 325877 165548 325924 165552
rect 325988 165550 326034 165610
rect 343174 165550 343220 165610
rect 343284 165608 343331 165612
rect 343326 165552 343331 165608
rect 325988 165548 325994 165550
rect 343214 165548 343220 165550
rect 343284 165548 343331 165552
rect 343398 165548 343404 165612
rect 343468 165610 343515 165612
rect 397453 165610 397519 165613
rect 398230 165610 398236 165612
rect 343468 165608 343560 165610
rect 343510 165552 343560 165608
rect 343468 165550 343560 165552
rect 397453 165608 398236 165610
rect 397453 165552 397458 165608
rect 397514 165552 398236 165608
rect 397453 165550 398236 165552
rect 343468 165548 343515 165550
rect 320909 165547 320975 165548
rect 325877 165547 325943 165548
rect 343265 165547 343331 165548
rect 343449 165547 343515 165548
rect 397453 165547 397519 165550
rect 398230 165548 398236 165550
rect 398300 165548 398306 165612
rect 401593 165610 401659 165613
rect 401726 165610 401732 165612
rect 401593 165608 401732 165610
rect 401593 165552 401598 165608
rect 401654 165552 401732 165608
rect 401593 165550 401732 165552
rect 401593 165547 401659 165550
rect 401726 165548 401732 165550
rect 401796 165548 401802 165612
rect 404353 165610 404419 165613
rect 405406 165610 405412 165612
rect 404353 165608 405412 165610
rect 404353 165552 404358 165608
rect 404414 165552 405412 165608
rect 404353 165550 405412 165552
rect 404353 165547 404419 165550
rect 405406 165548 405412 165550
rect 405476 165548 405482 165612
rect 407113 165610 407179 165613
rect 408166 165610 408172 165612
rect 407113 165608 408172 165610
rect 407113 165552 407118 165608
rect 407174 165552 408172 165608
rect 407113 165550 408172 165552
rect 407113 165547 407179 165550
rect 408166 165548 408172 165550
rect 408236 165548 408242 165612
rect 415485 165610 415551 165613
rect 416037 165612 416103 165613
rect 415894 165610 415900 165612
rect 415485 165608 415900 165610
rect 415485 165552 415490 165608
rect 415546 165552 415900 165608
rect 415485 165550 415900 165552
rect 415485 165547 415551 165550
rect 415894 165548 415900 165550
rect 415964 165548 415970 165612
rect 416037 165608 416084 165612
rect 416148 165610 416154 165612
rect 418705 165610 418771 165613
rect 419390 165610 419396 165612
rect 416037 165552 416042 165608
rect 416037 165548 416084 165552
rect 416148 165550 416194 165610
rect 418705 165608 419396 165610
rect 418705 165552 418710 165608
rect 418766 165552 419396 165608
rect 418705 165550 419396 165552
rect 416148 165548 416154 165550
rect 416037 165547 416103 165548
rect 418705 165547 418771 165550
rect 419390 165548 419396 165550
rect 419460 165548 419466 165612
rect 423673 165610 423739 165613
rect 423806 165610 423812 165612
rect 423673 165608 423812 165610
rect 423673 165552 423678 165608
rect 423734 165552 423812 165608
rect 423673 165550 423812 165552
rect 423673 165547 423739 165550
rect 423806 165548 423812 165550
rect 423876 165548 423882 165612
rect 426525 165610 426591 165613
rect 429653 165612 429719 165613
rect 427486 165610 427492 165612
rect 426525 165608 427492 165610
rect 426525 165552 426530 165608
rect 426586 165552 427492 165608
rect 426525 165550 427492 165552
rect 426525 165547 426591 165550
rect 427486 165548 427492 165550
rect 427556 165548 427562 165612
rect 429653 165608 429700 165612
rect 429764 165610 429770 165612
rect 435081 165610 435147 165613
rect 435909 165612 435975 165613
rect 437933 165612 437999 165613
rect 438485 165612 438551 165613
rect 435766 165610 435772 165612
rect 429653 165552 429658 165608
rect 429653 165548 429700 165552
rect 429764 165550 429810 165610
rect 435081 165608 435772 165610
rect 435081 165552 435086 165608
rect 435142 165552 435772 165608
rect 435081 165550 435772 165552
rect 429764 165548 429770 165550
rect 429653 165547 429719 165548
rect 435081 165547 435147 165550
rect 435766 165548 435772 165550
rect 435836 165548 435842 165612
rect 435909 165608 435956 165612
rect 436020 165610 436026 165612
rect 435909 165552 435914 165608
rect 435909 165548 435956 165552
rect 436020 165550 436066 165610
rect 437933 165608 437980 165612
rect 438044 165610 438050 165612
rect 437933 165552 437938 165608
rect 436020 165548 436026 165550
rect 437933 165548 437980 165552
rect 438044 165550 438090 165610
rect 438485 165608 438532 165612
rect 438596 165610 438602 165612
rect 438485 165552 438490 165608
rect 438044 165548 438050 165550
rect 438485 165548 438532 165552
rect 438596 165550 438642 165610
rect 438596 165548 438602 165550
rect 439262 165548 439268 165612
rect 439332 165610 439338 165612
rect 440141 165610 440207 165613
rect 439332 165608 440207 165610
rect 439332 165552 440146 165608
rect 440202 165552 440207 165608
rect 439332 165550 440207 165552
rect 439332 165548 439338 165550
rect 435909 165547 435975 165548
rect 437933 165547 437999 165548
rect 438485 165547 438551 165548
rect 440141 165547 440207 165550
rect 440877 165612 440943 165613
rect 443453 165612 443519 165613
rect 445845 165612 445911 165613
rect 440877 165608 440924 165612
rect 440988 165610 440994 165612
rect 440877 165552 440882 165608
rect 440877 165548 440924 165552
rect 440988 165550 441034 165610
rect 443453 165608 443500 165612
rect 443564 165610 443570 165612
rect 443453 165552 443458 165608
rect 440988 165548 440994 165550
rect 443453 165548 443500 165552
rect 443564 165550 443610 165610
rect 445845 165608 445892 165612
rect 445956 165610 445962 165612
rect 447317 165610 447383 165613
rect 448278 165610 448284 165612
rect 445845 165552 445850 165608
rect 443564 165548 443570 165550
rect 445845 165548 445892 165552
rect 445956 165550 446002 165610
rect 447317 165608 448284 165610
rect 447317 165552 447322 165608
rect 447378 165552 448284 165608
rect 447317 165550 448284 165552
rect 445956 165548 445962 165550
rect 440877 165547 440943 165548
rect 443453 165547 443519 165548
rect 445845 165547 445911 165548
rect 447317 165547 447383 165550
rect 448278 165548 448284 165550
rect 448348 165548 448354 165612
rect 449893 165610 449959 165613
rect 451038 165610 451044 165612
rect 449893 165608 451044 165610
rect 449893 165552 449898 165608
rect 449954 165552 451044 165608
rect 449893 165550 451044 165552
rect 449893 165547 449959 165550
rect 451038 165548 451044 165550
rect 451108 165548 451114 165612
rect 452653 165610 452719 165613
rect 453430 165610 453436 165612
rect 452653 165608 453436 165610
rect 452653 165552 452658 165608
rect 452714 165552 453436 165608
rect 452653 165550 453436 165552
rect 452653 165547 452719 165550
rect 453430 165548 453436 165550
rect 453500 165548 453506 165612
rect 455413 165610 455479 165613
rect 458357 165612 458423 165613
rect 503345 165612 503411 165613
rect 455822 165610 455828 165612
rect 455413 165608 455828 165610
rect 455413 165552 455418 165608
rect 455474 165552 455828 165608
rect 455413 165550 455828 165552
rect 455413 165547 455479 165550
rect 455822 165548 455828 165550
rect 455892 165548 455898 165612
rect 458357 165608 458404 165612
rect 458468 165610 458474 165612
rect 458357 165552 458362 165608
rect 458357 165548 458404 165552
rect 458468 165550 458514 165610
rect 458468 165548 458474 165550
rect 503294 165548 503300 165612
rect 503364 165610 503411 165612
rect 503364 165608 503456 165610
rect 503406 165552 503456 165608
rect 503364 165550 503456 165552
rect 503364 165548 503411 165550
rect 458357 165547 458423 165548
rect 503345 165547 503411 165548
rect 49233 165474 49299 165477
rect 158478 165474 158484 165476
rect 49233 165472 158484 165474
rect 49233 165416 49238 165472
rect 49294 165416 158484 165472
rect 49233 165414 158484 165416
rect 49233 165411 49299 165414
rect 158478 165412 158484 165414
rect 158548 165412 158554 165476
rect 166022 165412 166028 165476
rect 166092 165474 166098 165476
rect 198774 165474 198780 165476
rect 166092 165414 198780 165474
rect 166092 165412 166098 165414
rect 198774 165412 198780 165414
rect 198844 165412 198850 165476
rect 205214 165412 205220 165476
rect 205284 165474 205290 165476
rect 315798 165474 315804 165476
rect 205284 165414 315804 165474
rect 205284 165412 205290 165414
rect 315798 165412 315804 165414
rect 315868 165412 315874 165476
rect 378777 165474 378843 165477
rect 468518 165474 468524 165476
rect 378777 165472 468524 165474
rect 378777 165416 378782 165472
rect 378838 165416 468524 165472
rect 378777 165414 468524 165416
rect 378777 165411 378843 165414
rect 468518 165412 468524 165414
rect 468588 165412 468594 165476
rect 49325 165338 49391 165341
rect 155902 165338 155908 165340
rect 49325 165336 155908 165338
rect 49325 165280 49330 165336
rect 49386 165280 155908 165336
rect 49325 165278 155908 165280
rect 49325 165275 49391 165278
rect 155902 165276 155908 165278
rect 155972 165276 155978 165340
rect 206318 165276 206324 165340
rect 206388 165338 206394 165340
rect 311014 165338 311020 165340
rect 206388 165278 311020 165338
rect 206388 165276 206394 165278
rect 311014 165276 311020 165278
rect 311084 165276 311090 165340
rect 376017 165338 376083 165341
rect 465942 165338 465948 165340
rect 376017 165336 465948 165338
rect 376017 165280 376022 165336
rect 376078 165280 465948 165336
rect 376017 165278 465948 165280
rect 376017 165275 376083 165278
rect 465942 165276 465948 165278
rect 466012 165276 466018 165340
rect 49509 165202 49575 165205
rect 160870 165202 160876 165204
rect 49509 165200 160876 165202
rect 49509 165144 49514 165200
rect 49570 165144 160876 165200
rect 49509 165142 160876 165144
rect 49509 165139 49575 165142
rect 160870 165140 160876 165142
rect 160940 165140 160946 165204
rect 208158 165140 208164 165204
rect 208228 165202 208234 165204
rect 263726 165202 263732 165204
rect 208228 165142 263732 165202
rect 208228 165140 208234 165142
rect 263726 165140 263732 165142
rect 263796 165140 263802 165204
rect 264973 165202 265039 165205
rect 265198 165202 265204 165204
rect 264973 165200 265204 165202
rect 264973 165144 264978 165200
rect 265034 165144 265204 165200
rect 264973 165142 265204 165144
rect 264973 165139 265039 165142
rect 265198 165140 265204 165142
rect 265268 165140 265274 165204
rect 267733 165202 267799 165205
rect 268326 165202 268332 165204
rect 267733 165200 268332 165202
rect 267733 165144 267738 165200
rect 267794 165144 268332 165200
rect 267733 165142 268332 165144
rect 267733 165139 267799 165142
rect 268326 165140 268332 165142
rect 268396 165140 268402 165204
rect 271873 165202 271939 165205
rect 272190 165202 272196 165204
rect 271873 165200 272196 165202
rect 271873 165144 271878 165200
rect 271934 165144 272196 165200
rect 271873 165142 272196 165144
rect 271873 165139 271939 165142
rect 272190 165140 272196 165142
rect 272260 165140 272266 165204
rect 274817 165202 274883 165205
rect 276013 165204 276079 165205
rect 275686 165202 275692 165204
rect 274817 165200 275692 165202
rect 274817 165144 274822 165200
rect 274878 165144 275692 165200
rect 274817 165142 275692 165144
rect 274817 165139 274883 165142
rect 275686 165140 275692 165142
rect 275756 165140 275762 165204
rect 276013 165202 276060 165204
rect 275968 165200 276060 165202
rect 275968 165144 276018 165200
rect 275968 165142 276060 165144
rect 276013 165140 276060 165142
rect 276124 165140 276130 165204
rect 279182 165140 279188 165204
rect 279252 165202 279258 165204
rect 280061 165202 280127 165205
rect 279252 165200 280127 165202
rect 279252 165144 280066 165200
rect 280122 165144 280127 165200
rect 279252 165142 280127 165144
rect 279252 165140 279258 165142
rect 276013 165139 276079 165140
rect 280061 165139 280127 165142
rect 374862 165140 374868 165204
rect 374932 165202 374938 165204
rect 463550 165202 463556 165204
rect 374932 165142 463556 165202
rect 374932 165140 374938 165142
rect 463550 165140 463556 165142
rect 463620 165140 463626 165204
rect 118877 165066 118943 165069
rect 273437 165068 273503 165069
rect 432229 165068 432295 165069
rect 119102 165066 119108 165068
rect 118877 165064 119108 165066
rect 118877 165008 118882 165064
rect 118938 165008 119108 165064
rect 118877 165006 119108 165008
rect 118877 165003 118943 165006
rect 119102 165004 119108 165006
rect 119172 165004 119178 165068
rect 273437 165066 273484 165068
rect 273392 165064 273484 165066
rect 273392 165008 273442 165064
rect 273392 165006 273484 165008
rect 273437 165004 273484 165006
rect 273548 165004 273554 165068
rect 379462 165004 379468 165068
rect 379532 165066 379538 165068
rect 426014 165066 426020 165068
rect 379532 165006 426020 165066
rect 379532 165004 379538 165006
rect 426014 165004 426020 165006
rect 426084 165004 426090 165068
rect 432229 165064 432276 165068
rect 432340 165066 432346 165068
rect 432229 165008 432234 165064
rect 432229 165004 432276 165008
rect 432340 165006 432386 165066
rect 432340 165004 432346 165006
rect 273437 165003 273503 165004
rect 432229 165003 432295 165004
rect 114461 164932 114527 164933
rect 114461 164928 114508 164932
rect 114572 164930 114578 164932
rect 247033 164930 247099 164933
rect 248270 164930 248276 164932
rect 114461 164872 114466 164928
rect 114461 164868 114508 164872
rect 114572 164870 114618 164930
rect 247033 164928 248276 164930
rect 247033 164872 247038 164928
rect 247094 164872 248276 164928
rect 247033 164870 248276 164872
rect 114572 164868 114578 164870
rect 114461 164867 114527 164868
rect 247033 164867 247099 164870
rect 248270 164868 248276 164870
rect 248340 164868 248346 164932
rect 249793 164930 249859 164933
rect 250662 164930 250668 164932
rect 249793 164928 250668 164930
rect 249793 164872 249798 164928
rect 249854 164872 250668 164928
rect 249793 164870 250668 164872
rect 249793 164867 249859 164870
rect 250662 164868 250668 164870
rect 250732 164868 250738 164932
rect 252553 164930 252619 164933
rect 253606 164930 253612 164932
rect 252553 164928 253612 164930
rect 252553 164872 252558 164928
rect 252614 164872 253612 164928
rect 252553 164870 253612 164872
rect 252553 164867 252619 164870
rect 253606 164868 253612 164870
rect 253676 164868 253682 164932
rect 258073 164930 258139 164933
rect 258390 164930 258396 164932
rect 258073 164928 258396 164930
rect 258073 164872 258078 164928
rect 258134 164872 258396 164928
rect 258073 164870 258396 164872
rect 258073 164867 258139 164870
rect 258390 164868 258396 164870
rect 258460 164868 258466 164932
rect 412633 164930 412699 164933
rect 413686 164930 413692 164932
rect 412633 164928 413692 164930
rect 412633 164872 412638 164928
rect 412694 164872 413692 164928
rect 412633 164870 413692 164872
rect 412633 164867 412699 164870
rect 413686 164868 413692 164870
rect 413756 164868 413762 164932
rect 436185 164930 436251 164933
rect 436870 164930 436876 164932
rect 436185 164928 436876 164930
rect 436185 164872 436190 164928
rect 436246 164872 436876 164928
rect 436185 164870 436876 164872
rect 436185 164867 436251 164870
rect 436870 164868 436876 164870
rect 436940 164868 436946 164932
rect 88333 164796 88399 164797
rect 88333 164794 88380 164796
rect 88288 164792 88380 164794
rect 88288 164736 88338 164792
rect 88288 164734 88380 164736
rect 88333 164732 88380 164734
rect 88444 164732 88450 164796
rect 89989 164794 90055 164797
rect 90766 164794 90772 164796
rect 89989 164792 90772 164794
rect 89989 164736 89994 164792
rect 90050 164736 90772 164792
rect 89989 164734 90772 164736
rect 88333 164731 88399 164732
rect 89989 164731 90055 164734
rect 90766 164732 90772 164734
rect 90836 164732 90842 164796
rect 200982 164732 200988 164796
rect 201052 164794 201058 164796
rect 323342 164794 323348 164796
rect 201052 164734 323348 164794
rect 201052 164732 201058 164734
rect 323342 164732 323348 164734
rect 323412 164732 323418 164796
rect 409873 164794 409939 164797
rect 410742 164794 410748 164796
rect 409873 164792 410748 164794
rect 409873 164736 409878 164792
rect 409934 164736 410748 164792
rect 409873 164734 410748 164736
rect 409873 164731 409939 164734
rect 410742 164732 410748 164734
rect 410812 164732 410818 164796
rect 112069 164660 112135 164661
rect 115749 164660 115815 164661
rect 112069 164656 112116 164660
rect 112180 164658 112186 164660
rect 112069 164600 112074 164656
rect 112069 164596 112116 164600
rect 112180 164598 112226 164658
rect 115749 164656 115796 164660
rect 115860 164658 115866 164660
rect 369301 164658 369367 164661
rect 460974 164658 460980 164660
rect 115749 164600 115754 164656
rect 112180 164596 112186 164598
rect 115749 164596 115796 164600
rect 115860 164598 115906 164658
rect 369301 164656 460980 164658
rect 369301 164600 369306 164656
rect 369362 164600 460980 164656
rect 369301 164598 460980 164600
rect 115860 164596 115866 164598
rect 112069 164595 112135 164596
rect 115749 164595 115815 164596
rect 369301 164595 369367 164598
rect 460974 164596 460980 164598
rect 461044 164596 461050 164660
rect 96613 164522 96679 164525
rect 97022 164522 97028 164524
rect 96613 164520 97028 164522
rect 96613 164464 96618 164520
rect 96674 164464 97028 164520
rect 96613 164462 97028 164464
rect 96613 164459 96679 164462
rect 97022 164460 97028 164462
rect 97092 164460 97098 164524
rect 113214 164460 113220 164524
rect 113284 164522 113290 164524
rect 114645 164522 114711 164525
rect 113284 164520 114711 164522
rect 113284 164464 114650 164520
rect 114706 164464 114711 164520
rect 113284 164462 114711 164464
rect 113284 164460 113290 164462
rect 114645 164459 114711 164462
rect 420913 164522 420979 164525
rect 421782 164522 421788 164524
rect 420913 164520 421788 164522
rect 420913 164464 420918 164520
rect 420974 164464 421788 164520
rect 420913 164462 421788 164464
rect 420913 164459 420979 164462
rect 421782 164460 421788 164462
rect 421852 164460 421858 164524
rect 430573 164522 430639 164525
rect 431166 164522 431172 164524
rect 430573 164520 431172 164522
rect 430573 164464 430578 164520
rect 430634 164464 431172 164520
rect 430573 164462 431172 164464
rect 430573 164459 430639 164462
rect 431166 164460 431172 164462
rect 431236 164460 431242 164524
rect 75913 164386 75979 164389
rect 77150 164386 77156 164388
rect 75913 164384 77156 164386
rect 75913 164328 75918 164384
rect 75974 164328 77156 164384
rect 75913 164326 77156 164328
rect 75913 164323 75979 164326
rect 77150 164324 77156 164326
rect 77220 164324 77226 164388
rect 100753 164386 100819 164389
rect 101806 164386 101812 164388
rect 100753 164384 101812 164386
rect 100753 164328 100758 164384
rect 100814 164328 101812 164384
rect 100753 164326 101812 164328
rect 100753 164323 100819 164326
rect 101806 164324 101812 164326
rect 101876 164324 101882 164388
rect 103513 164386 103579 164389
rect 103830 164386 103836 164388
rect 103513 164384 103836 164386
rect 103513 164328 103518 164384
rect 103574 164328 103836 164384
rect 103513 164326 103836 164328
rect 103513 164323 103579 164326
rect 103830 164324 103836 164326
rect 103900 164324 103906 164388
rect 244273 164386 244339 164389
rect 244406 164386 244412 164388
rect 244273 164384 244412 164386
rect 244273 164328 244278 164384
rect 244334 164328 244412 164384
rect 244273 164326 244412 164328
rect 244273 164323 244339 164326
rect 244406 164324 244412 164326
rect 244476 164324 244482 164388
rect 251265 164386 251331 164389
rect 252318 164386 252324 164388
rect 251265 164384 252324 164386
rect 251265 164328 251270 164384
rect 251326 164328 252324 164384
rect 251265 164326 252324 164328
rect 251265 164323 251331 164326
rect 252318 164324 252324 164326
rect 252388 164324 252394 164388
rect 259545 164386 259611 164389
rect 260598 164386 260604 164388
rect 259545 164384 260604 164386
rect 259545 164328 259550 164384
rect 259606 164328 260604 164384
rect 259545 164326 260604 164328
rect 259545 164323 259611 164326
rect 260598 164324 260604 164326
rect 260668 164324 260674 164388
rect 266486 164324 266492 164388
rect 266556 164386 266562 164388
rect 267641 164386 267707 164389
rect 266556 164384 267707 164386
rect 266556 164328 267646 164384
rect 267702 164328 267707 164384
rect 266556 164326 267707 164328
rect 266556 164324 266562 164326
rect 267641 164323 267707 164326
rect 273805 164386 273871 164389
rect 274398 164386 274404 164388
rect 273805 164384 274404 164386
rect 273805 164328 273810 164384
rect 273866 164328 274404 164384
rect 273805 164326 274404 164328
rect 273805 164323 273871 164326
rect 274398 164324 274404 164326
rect 274468 164324 274474 164388
rect 396165 164386 396231 164389
rect 397126 164386 397132 164388
rect 396165 164384 397132 164386
rect 396165 164328 396170 164384
rect 396226 164328 397132 164384
rect 396165 164326 397132 164328
rect 396165 164323 396231 164326
rect 397126 164324 397132 164326
rect 397196 164324 397202 164388
rect 403065 164386 403131 164389
rect 404118 164386 404124 164388
rect 403065 164384 404124 164386
rect 403065 164328 403070 164384
rect 403126 164328 404124 164384
rect 403065 164326 404124 164328
rect 403065 164323 403131 164326
rect 404118 164324 404124 164326
rect 404188 164324 404194 164388
rect 411345 164386 411411 164389
rect 412398 164386 412404 164388
rect 411345 164384 412404 164386
rect 411345 164328 411350 164384
rect 411406 164328 412404 164384
rect 411345 164326 412404 164328
rect 411345 164323 411411 164326
rect 412398 164324 412404 164326
rect 412468 164324 412474 164388
rect 76005 164252 76071 164253
rect 76005 164248 76052 164252
rect 76116 164250 76122 164252
rect 77293 164250 77359 164253
rect 78254 164250 78260 164252
rect 76005 164192 76010 164248
rect 76005 164188 76052 164192
rect 76116 164190 76162 164250
rect 77293 164248 78260 164250
rect 77293 164192 77298 164248
rect 77354 164192 78260 164248
rect 77293 164190 78260 164192
rect 76116 164188 76122 164190
rect 76005 164187 76071 164188
rect 77293 164187 77359 164190
rect 78254 164188 78260 164190
rect 78324 164188 78330 164252
rect 78673 164250 78739 164253
rect 79542 164250 79548 164252
rect 78673 164248 79548 164250
rect 78673 164192 78678 164248
rect 78734 164192 79548 164248
rect 78673 164190 79548 164192
rect 78673 164187 78739 164190
rect 79542 164188 79548 164190
rect 79612 164188 79618 164252
rect 80053 164250 80119 164253
rect 80462 164250 80468 164252
rect 80053 164248 80468 164250
rect 80053 164192 80058 164248
rect 80114 164192 80468 164248
rect 80053 164190 80468 164192
rect 80053 164187 80119 164190
rect 80462 164188 80468 164190
rect 80532 164188 80538 164252
rect 82813 164250 82879 164253
rect 83038 164250 83044 164252
rect 82813 164248 83044 164250
rect 82813 164192 82818 164248
rect 82874 164192 83044 164248
rect 82813 164190 83044 164192
rect 82813 164187 82879 164190
rect 83038 164188 83044 164190
rect 83108 164188 83114 164252
rect 84142 164188 84148 164252
rect 84212 164250 84218 164252
rect 84285 164250 84351 164253
rect 84212 164248 84351 164250
rect 84212 164192 84290 164248
rect 84346 164192 84351 164248
rect 84212 164190 84351 164192
rect 84212 164188 84218 164190
rect 84285 164187 84351 164190
rect 85573 164250 85639 164253
rect 86534 164250 86540 164252
rect 85573 164248 86540 164250
rect 85573 164192 85578 164248
rect 85634 164192 86540 164248
rect 85573 164190 86540 164192
rect 85573 164187 85639 164190
rect 86534 164188 86540 164190
rect 86604 164188 86610 164252
rect 86953 164250 87019 164253
rect 87638 164250 87644 164252
rect 86953 164248 87644 164250
rect 86953 164192 86958 164248
rect 87014 164192 87644 164248
rect 86953 164190 87644 164192
rect 86953 164187 87019 164190
rect 87638 164188 87644 164190
rect 87708 164188 87714 164252
rect 88425 164250 88491 164253
rect 88742 164250 88748 164252
rect 88425 164248 88748 164250
rect 88425 164192 88430 164248
rect 88486 164192 88748 164248
rect 88425 164190 88748 164192
rect 88425 164187 88491 164190
rect 88742 164188 88748 164190
rect 88812 164188 88818 164252
rect 89805 164250 89871 164253
rect 90030 164250 90036 164252
rect 89805 164248 90036 164250
rect 89805 164192 89810 164248
rect 89866 164192 90036 164248
rect 89805 164190 90036 164192
rect 89805 164187 89871 164190
rect 90030 164188 90036 164190
rect 90100 164188 90106 164252
rect 91093 164250 91159 164253
rect 91318 164250 91324 164252
rect 91093 164248 91324 164250
rect 91093 164192 91098 164248
rect 91154 164192 91324 164248
rect 91093 164190 91324 164192
rect 91093 164187 91159 164190
rect 91318 164188 91324 164190
rect 91388 164188 91394 164252
rect 92473 164250 92539 164253
rect 93342 164250 93348 164252
rect 92473 164248 93348 164250
rect 92473 164192 92478 164248
rect 92534 164192 93348 164248
rect 92473 164190 93348 164192
rect 92473 164187 92539 164190
rect 93342 164188 93348 164190
rect 93412 164188 93418 164252
rect 93853 164250 93919 164253
rect 94446 164250 94452 164252
rect 93853 164248 94452 164250
rect 93853 164192 93858 164248
rect 93914 164192 94452 164248
rect 93853 164190 94452 164192
rect 93853 164187 93919 164190
rect 94446 164188 94452 164190
rect 94516 164188 94522 164252
rect 97993 164250 98059 164253
rect 100753 164252 100819 164253
rect 98126 164250 98132 164252
rect 97993 164248 98132 164250
rect 97993 164192 97998 164248
rect 98054 164192 98132 164248
rect 97993 164190 98132 164192
rect 97993 164187 98059 164190
rect 98126 164188 98132 164190
rect 98196 164188 98202 164252
rect 100702 164250 100708 164252
rect 100662 164190 100708 164250
rect 100772 164248 100819 164252
rect 100814 164192 100819 164248
rect 100702 164188 100708 164190
rect 100772 164188 100819 164192
rect 100753 164187 100819 164188
rect 102133 164250 102199 164253
rect 102726 164250 102732 164252
rect 102133 164248 102732 164250
rect 102133 164192 102138 164248
rect 102194 164192 102732 164248
rect 102133 164190 102732 164192
rect 102133 164187 102199 164190
rect 102726 164188 102732 164190
rect 102796 164188 102802 164252
rect 105302 164188 105308 164252
rect 105372 164250 105378 164252
rect 106181 164250 106247 164253
rect 105372 164248 106247 164250
rect 105372 164192 106186 164248
rect 106242 164192 106247 164248
rect 105372 164190 106247 164192
rect 105372 164188 105378 164190
rect 106181 164187 106247 164190
rect 106365 164252 106431 164253
rect 107561 164252 107627 164253
rect 106365 164248 106412 164252
rect 106476 164250 106482 164252
rect 107510 164250 107516 164252
rect 106365 164192 106370 164248
rect 106365 164188 106412 164192
rect 106476 164190 106522 164250
rect 107470 164190 107516 164250
rect 107580 164248 107627 164252
rect 108614 164250 108620 164252
rect 107622 164192 107627 164248
rect 106476 164188 106482 164190
rect 107510 164188 107516 164190
rect 107580 164188 107627 164192
rect 106365 164187 106431 164188
rect 107561 164187 107627 164188
rect 107702 164190 108620 164250
rect 107702 164117 107762 164190
rect 108614 164188 108620 164190
rect 108684 164188 108690 164252
rect 235993 164250 236059 164253
rect 237046 164250 237052 164252
rect 235993 164248 237052 164250
rect 235993 164192 235998 164248
rect 236054 164192 237052 164248
rect 235993 164190 237052 164192
rect 235993 164187 236059 164190
rect 237046 164188 237052 164190
rect 237116 164188 237122 164252
rect 237373 164250 237439 164253
rect 238150 164250 238156 164252
rect 237373 164248 238156 164250
rect 237373 164192 237378 164248
rect 237434 164192 238156 164248
rect 237373 164190 238156 164192
rect 237373 164187 237439 164190
rect 238150 164188 238156 164190
rect 238220 164188 238226 164252
rect 240133 164250 240199 164253
rect 240542 164250 240548 164252
rect 240133 164248 240548 164250
rect 240133 164192 240138 164248
rect 240194 164192 240548 164248
rect 240133 164190 240548 164192
rect 240133 164187 240199 164190
rect 240542 164188 240548 164190
rect 240612 164188 240618 164252
rect 241513 164250 241579 164253
rect 241646 164250 241652 164252
rect 241513 164248 241652 164250
rect 241513 164192 241518 164248
rect 241574 164192 241652 164248
rect 241513 164190 241652 164192
rect 241513 164187 241579 164190
rect 241646 164188 241652 164190
rect 241716 164188 241722 164252
rect 244365 164250 244431 164253
rect 245326 164250 245332 164252
rect 244365 164248 245332 164250
rect 244365 164192 244370 164248
rect 244426 164192 245332 164248
rect 244365 164190 245332 164192
rect 244365 164187 244431 164190
rect 245326 164188 245332 164190
rect 245396 164188 245402 164252
rect 245653 164250 245719 164253
rect 246430 164250 246436 164252
rect 245653 164248 246436 164250
rect 245653 164192 245658 164248
rect 245714 164192 246436 164248
rect 245653 164190 246436 164192
rect 245653 164187 245719 164190
rect 246430 164188 246436 164190
rect 246500 164188 246506 164252
rect 248413 164250 248479 164253
rect 248638 164250 248644 164252
rect 248413 164248 248644 164250
rect 248413 164192 248418 164248
rect 248474 164192 248644 164248
rect 248413 164190 248644 164192
rect 248413 164187 248479 164190
rect 248638 164188 248644 164190
rect 248708 164188 248714 164252
rect 249885 164250 249951 164253
rect 251173 164252 251239 164253
rect 250110 164250 250116 164252
rect 249885 164248 250116 164250
rect 249885 164192 249890 164248
rect 249946 164192 250116 164248
rect 249885 164190 250116 164192
rect 249885 164187 249951 164190
rect 250110 164188 250116 164190
rect 250180 164188 250186 164252
rect 251173 164250 251220 164252
rect 251128 164248 251220 164250
rect 251128 164192 251178 164248
rect 251128 164190 251220 164192
rect 251173 164188 251220 164190
rect 251284 164188 251290 164252
rect 252645 164250 252711 164253
rect 253422 164250 253428 164252
rect 252645 164248 253428 164250
rect 252645 164192 252650 164248
rect 252706 164192 253428 164248
rect 252645 164190 253428 164192
rect 251173 164187 251239 164188
rect 252645 164187 252711 164190
rect 253422 164188 253428 164190
rect 253492 164188 253498 164252
rect 253933 164250 253999 164253
rect 254526 164250 254532 164252
rect 253933 164248 254532 164250
rect 253933 164192 253938 164248
rect 253994 164192 254532 164248
rect 253933 164190 254532 164192
rect 253933 164187 253999 164190
rect 254526 164188 254532 164190
rect 254596 164188 254602 164252
rect 255405 164250 255471 164253
rect 255814 164250 255820 164252
rect 255405 164248 255820 164250
rect 255405 164192 255410 164248
rect 255466 164192 255820 164248
rect 255405 164190 255820 164192
rect 255405 164187 255471 164190
rect 255814 164188 255820 164190
rect 255884 164188 255890 164252
rect 256693 164250 256759 164253
rect 259453 164252 259519 164253
rect 256918 164250 256924 164252
rect 256693 164248 256924 164250
rect 256693 164192 256698 164248
rect 256754 164192 256924 164248
rect 256693 164190 256924 164192
rect 256693 164187 256759 164190
rect 256918 164188 256924 164190
rect 256988 164188 256994 164252
rect 259453 164250 259500 164252
rect 259408 164248 259500 164250
rect 259408 164192 259458 164248
rect 259408 164190 259500 164192
rect 259453 164188 259500 164190
rect 259564 164188 259570 164252
rect 262806 164188 262812 164252
rect 262876 164250 262882 164252
rect 263501 164250 263567 164253
rect 262876 164248 263567 164250
rect 262876 164192 263506 164248
rect 263562 164192 263567 164248
rect 262876 164190 263567 164192
rect 262876 164188 262882 164190
rect 259453 164187 259519 164188
rect 263501 164187 263567 164190
rect 263777 164250 263843 164253
rect 263910 164250 263916 164252
rect 263777 164248 263916 164250
rect 263777 164192 263782 164248
rect 263838 164192 263916 164248
rect 263777 164190 263916 164192
rect 263777 164187 263843 164190
rect 263910 164188 263916 164190
rect 263980 164188 263986 164252
rect 266353 164250 266419 164253
rect 267590 164250 267596 164252
rect 266353 164248 267596 164250
rect 266353 164192 266358 164248
rect 266414 164192 267596 164248
rect 266353 164190 267596 164192
rect 266353 164187 266419 164190
rect 267590 164188 267596 164190
rect 267660 164188 267666 164252
rect 267733 164250 267799 164253
rect 268694 164250 268700 164252
rect 267733 164248 268700 164250
rect 267733 164192 267738 164248
rect 267794 164192 268700 164248
rect 267733 164190 268700 164192
rect 267733 164187 267799 164190
rect 268694 164188 268700 164190
rect 268764 164188 268770 164252
rect 269113 164250 269179 164253
rect 269798 164250 269804 164252
rect 269113 164248 269804 164250
rect 269113 164192 269118 164248
rect 269174 164192 269804 164248
rect 269113 164190 269804 164192
rect 269113 164187 269179 164190
rect 269798 164188 269804 164190
rect 269868 164188 269874 164252
rect 270493 164250 270559 164253
rect 271270 164250 271276 164252
rect 270493 164248 271276 164250
rect 270493 164192 270498 164248
rect 270554 164192 271276 164248
rect 270493 164190 271276 164192
rect 270493 164187 270559 164190
rect 271270 164188 271276 164190
rect 271340 164188 271346 164252
rect 273294 164188 273300 164252
rect 273364 164250 273370 164252
rect 274541 164250 274607 164253
rect 273364 164248 274607 164250
rect 273364 164192 274546 164248
rect 274602 164192 274607 164248
rect 273364 164190 274607 164192
rect 273364 164188 273370 164190
rect 274541 164187 274607 164190
rect 276974 164188 276980 164252
rect 277044 164250 277050 164252
rect 277301 164250 277367 164253
rect 278037 164252 278103 164253
rect 396073 164252 396139 164253
rect 278037 164250 278084 164252
rect 277044 164248 277367 164250
rect 277044 164192 277306 164248
rect 277362 164192 277367 164248
rect 277044 164190 277367 164192
rect 277992 164248 278084 164250
rect 277992 164192 278042 164248
rect 277992 164190 278084 164192
rect 277044 164188 277050 164190
rect 277301 164187 277367 164190
rect 278037 164188 278084 164190
rect 278148 164188 278154 164252
rect 318374 164250 318380 164252
rect 315990 164190 318380 164250
rect 278037 164187 278103 164188
rect 57513 164116 57579 164117
rect 57462 164052 57468 164116
rect 57532 164114 57579 164116
rect 57532 164112 57624 164114
rect 57574 164056 57624 164112
rect 57532 164054 57624 164056
rect 107653 164112 107762 164117
rect 107653 164056 107658 164112
rect 107714 164056 107762 164112
rect 107653 164054 107762 164056
rect 57532 164052 57579 164054
rect 57513 164051 57579 164052
rect 107653 164051 107719 164054
rect 214598 164052 214604 164116
rect 214668 164114 214674 164116
rect 315990 164114 316050 164190
rect 318374 164188 318380 164190
rect 318444 164188 318450 164252
rect 396022 164250 396028 164252
rect 395982 164190 396028 164250
rect 396092 164248 396139 164252
rect 396134 164192 396139 164248
rect 396022 164188 396028 164190
rect 396092 164188 396139 164192
rect 396073 164187 396139 164188
rect 398833 164250 398899 164253
rect 399518 164250 399524 164252
rect 398833 164248 399524 164250
rect 398833 164192 398838 164248
rect 398894 164192 399524 164248
rect 398833 164190 399524 164192
rect 398833 164187 398899 164190
rect 399518 164188 399524 164190
rect 399588 164188 399594 164252
rect 400213 164250 400279 164253
rect 402973 164252 403039 164253
rect 400438 164250 400444 164252
rect 400213 164248 400444 164250
rect 400213 164192 400218 164248
rect 400274 164192 400444 164248
rect 400213 164190 400444 164192
rect 400213 164187 400279 164190
rect 400438 164188 400444 164190
rect 400508 164188 400514 164252
rect 402973 164250 403020 164252
rect 402928 164248 403020 164250
rect 402928 164192 402978 164248
rect 402928 164190 403020 164192
rect 402973 164188 403020 164190
rect 403084 164188 403090 164252
rect 405733 164250 405799 164253
rect 406510 164250 406516 164252
rect 405733 164248 406516 164250
rect 405733 164192 405738 164248
rect 405794 164192 406516 164248
rect 405733 164190 406516 164192
rect 402973 164187 403039 164188
rect 405733 164187 405799 164190
rect 406510 164188 406516 164190
rect 406580 164188 406586 164252
rect 407205 164250 407271 164253
rect 407614 164250 407620 164252
rect 407205 164248 407620 164250
rect 407205 164192 407210 164248
rect 407266 164192 407620 164248
rect 407205 164190 407620 164192
rect 407205 164187 407271 164190
rect 407614 164188 407620 164190
rect 407684 164188 407690 164252
rect 408493 164250 408559 164253
rect 409965 164252 410031 164253
rect 411253 164252 411319 164253
rect 408718 164250 408724 164252
rect 408493 164248 408724 164250
rect 408493 164192 408498 164248
rect 408554 164192 408724 164248
rect 408493 164190 408724 164192
rect 408493 164187 408559 164190
rect 408718 164188 408724 164190
rect 408788 164188 408794 164252
rect 409965 164250 410012 164252
rect 409920 164248 410012 164250
rect 409920 164192 409970 164248
rect 409920 164190 410012 164192
rect 409965 164188 410012 164190
rect 410076 164188 410082 164252
rect 411253 164250 411300 164252
rect 411208 164248 411300 164250
rect 411208 164192 411258 164248
rect 411208 164190 411300 164192
rect 411253 164188 411300 164190
rect 411364 164188 411370 164252
rect 412633 164250 412699 164253
rect 413318 164250 413324 164252
rect 412633 164248 413324 164250
rect 412633 164192 412638 164248
rect 412694 164192 413324 164248
rect 412633 164190 413324 164192
rect 409965 164187 410031 164188
rect 411253 164187 411319 164188
rect 412633 164187 412699 164190
rect 413318 164188 413324 164190
rect 413388 164188 413394 164252
rect 414013 164250 414079 164253
rect 414422 164250 414428 164252
rect 414013 164248 414428 164250
rect 414013 164192 414018 164248
rect 414074 164192 414428 164248
rect 414013 164190 414428 164192
rect 414013 164187 414079 164190
rect 414422 164188 414428 164190
rect 414492 164188 414498 164252
rect 416773 164250 416839 164253
rect 416998 164250 417004 164252
rect 416773 164248 417004 164250
rect 416773 164192 416778 164248
rect 416834 164192 417004 164248
rect 416773 164190 417004 164192
rect 416773 164187 416839 164190
rect 416998 164188 417004 164190
rect 417068 164188 417074 164252
rect 418153 164250 418219 164253
rect 418286 164250 418292 164252
rect 418153 164248 418292 164250
rect 418153 164192 418158 164248
rect 418214 164192 418292 164248
rect 418153 164190 418292 164192
rect 418153 164187 418219 164190
rect 418286 164188 418292 164190
rect 418356 164188 418362 164252
rect 419533 164250 419599 164253
rect 420678 164250 420684 164252
rect 419533 164248 420684 164250
rect 419533 164192 419538 164248
rect 419594 164192 420684 164248
rect 419533 164190 420684 164192
rect 419533 164187 419599 164190
rect 420678 164188 420684 164190
rect 420748 164188 420754 164252
rect 422293 164250 422359 164253
rect 422886 164250 422892 164252
rect 422293 164248 422892 164250
rect 422293 164192 422298 164248
rect 422354 164192 422892 164248
rect 422293 164190 422892 164192
rect 422293 164187 422359 164190
rect 422886 164188 422892 164190
rect 422956 164188 422962 164252
rect 425053 164250 425119 164253
rect 426433 164252 426499 164253
rect 425278 164250 425284 164252
rect 425053 164248 425284 164250
rect 425053 164192 425058 164248
rect 425114 164192 425284 164248
rect 425053 164190 425284 164192
rect 425053 164187 425119 164190
rect 425278 164188 425284 164190
rect 425348 164188 425354 164252
rect 426382 164188 426388 164252
rect 426452 164250 426499 164252
rect 426452 164248 426544 164250
rect 426494 164192 426544 164248
rect 426452 164190 426544 164192
rect 426452 164188 426499 164190
rect 428774 164188 428780 164252
rect 428844 164250 428850 164252
rect 429101 164250 429167 164253
rect 428844 164248 429167 164250
rect 428844 164192 429106 164248
rect 429162 164192 429167 164248
rect 428844 164190 429167 164192
rect 428844 164188 428850 164190
rect 426433 164187 426499 164188
rect 429101 164187 429167 164190
rect 433374 164188 433380 164252
rect 433444 164250 433450 164252
rect 434621 164250 434687 164253
rect 433444 164248 434687 164250
rect 433444 164192 434626 164248
rect 434682 164192 434687 164248
rect 433444 164190 434687 164192
rect 433444 164188 433450 164190
rect 434621 164187 434687 164190
rect 214668 164054 316050 164114
rect 214668 164052 214674 164054
rect 207974 163916 207980 163980
rect 208044 163978 208050 163980
rect 308213 163978 308279 163981
rect 208044 163976 308279 163978
rect 208044 163920 308218 163976
rect 308274 163920 308279 163976
rect 208044 163918 308279 163920
rect 208044 163916 208050 163918
rect 308213 163915 308279 163918
rect -960 162740 480 162980
rect 217174 162556 217180 162620
rect 217244 162618 217250 162620
rect 217317 162618 217383 162621
rect 217244 162616 217383 162618
rect 217244 162560 217322 162616
rect 217378 162560 217383 162616
rect 217244 162558 217383 162560
rect 217244 162556 217250 162558
rect 217317 162555 217383 162558
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect -960 149774 674 149834
rect -960 149698 480 149774
rect 614 149698 674 149774
rect -960 149684 674 149698
rect 246 149638 674 149684
rect 246 149154 306 149638
rect 360878 149154 360884 149156
rect 246 149094 360884 149154
rect 360878 149092 360884 149094
rect 360948 149092 360954 149156
rect 278037 149018 278103 149021
rect 278681 149018 278747 149021
rect 357433 149018 357499 149021
rect 278037 149016 357499 149018
rect 278037 148960 278042 149016
rect 278098 148960 278686 149016
rect 278742 148960 357438 149016
rect 357494 148960 357499 149016
rect 278037 148958 357499 148960
rect 278037 148955 278103 148958
rect 278681 148955 278747 148958
rect 357433 148955 357499 148958
rect 217358 148276 217364 148340
rect 217428 148338 217434 148340
rect 278681 148338 278747 148341
rect 217428 148336 278747 148338
rect 217428 148280 278686 148336
rect 278742 148280 278747 148336
rect 217428 148278 278747 148280
rect 217428 148276 217434 148278
rect 278681 148275 278747 148278
rect 377622 148276 377628 148340
rect 377692 148338 377698 148340
rect 440233 148338 440299 148341
rect 377692 148336 440299 148338
rect 377692 148280 440238 148336
rect 440294 148280 440299 148336
rect 377692 148278 440299 148280
rect 377692 148276 377698 148278
rect 440233 148275 440299 148278
rect 57646 147732 57652 147796
rect 57716 147794 57722 147796
rect 58709 147794 58775 147797
rect 57716 147792 58775 147794
rect 57716 147736 58714 147792
rect 58770 147736 58775 147792
rect 57716 147734 58775 147736
rect 57716 147732 57722 147734
rect 58709 147731 58775 147734
rect 56225 146298 56291 146301
rect 58801 146298 58867 146301
rect 102133 146298 102199 146301
rect 56225 146296 102199 146298
rect 56225 146240 56230 146296
rect 56286 146240 58806 146296
rect 58862 146240 102138 146296
rect 102194 146240 102199 146296
rect 56225 146238 102199 146240
rect 56225 146235 56291 146238
rect 58801 146235 58867 146238
rect 102133 146235 102199 146238
rect 214189 146298 214255 146301
rect 214925 146298 214991 146301
rect 269113 146298 269179 146301
rect 214189 146296 269179 146298
rect 214189 146240 214194 146296
rect 214250 146240 214930 146296
rect 214986 146240 269118 146296
rect 269174 146240 269179 146296
rect 214189 146238 269179 146240
rect 214189 146235 214255 146238
rect 214925 146235 214991 146238
rect 269113 146235 269179 146238
rect 377990 146236 377996 146300
rect 378060 146298 378066 146300
rect 378409 146298 378475 146301
rect 378060 146296 378475 146298
rect 378060 146240 378414 146296
rect 378470 146240 378475 146296
rect 378060 146238 378475 146240
rect 378060 146236 378066 146238
rect 378409 146235 378475 146238
rect 218605 146162 218671 146165
rect 267825 146162 267891 146165
rect 218605 146160 267891 146162
rect 218605 146104 218610 146160
rect 218666 146104 267830 146160
rect 267886 146104 267891 146160
rect 218605 146102 267891 146104
rect 218605 146099 218671 146102
rect 267825 146099 267891 146102
rect 372245 146162 372311 146165
rect 379462 146162 379468 146164
rect 372245 146160 379468 146162
rect 372245 146104 372250 146160
rect 372306 146104 379468 146160
rect 372245 146102 379468 146104
rect 372245 146099 372311 146102
rect 379462 146100 379468 146102
rect 379532 146100 379538 146164
rect 216581 146026 216647 146029
rect 263593 146026 263659 146029
rect 216581 146024 263659 146026
rect 216581 145968 216586 146024
rect 216642 145968 263598 146024
rect 263654 145968 263659 146024
rect 216581 145966 263659 145968
rect 216581 145963 216647 145966
rect 263593 145963 263659 145966
rect 378409 146026 378475 146029
rect 415485 146026 415551 146029
rect 378409 146024 415551 146026
rect 378409 145968 378414 146024
rect 378470 145968 415490 146024
rect 415546 145968 415551 146024
rect 378409 145966 415551 145968
rect 378409 145963 378475 145966
rect 415485 145963 415551 145966
rect 54477 145890 54543 145893
rect 58985 145890 59051 145893
rect 100753 145890 100819 145893
rect 54477 145888 100819 145890
rect 54477 145832 54482 145888
rect 54538 145832 58990 145888
rect 59046 145832 100758 145888
rect 100814 145832 100819 145888
rect 54477 145830 100819 145832
rect 54477 145827 54543 145830
rect 58985 145827 59051 145830
rect 100753 145827 100819 145830
rect 219893 145890 219959 145893
rect 220813 145890 220879 145893
rect 267733 145890 267799 145893
rect 219893 145888 267799 145890
rect 219893 145832 219898 145888
rect 219954 145832 220818 145888
rect 220874 145832 267738 145888
rect 267794 145832 267799 145888
rect 219893 145830 267799 145832
rect 219893 145827 219959 145830
rect 220813 145827 220879 145830
rect 267733 145827 267799 145830
rect 377949 145890 378015 145893
rect 423673 145890 423739 145893
rect 377949 145888 423739 145890
rect 377949 145832 377954 145888
rect 378010 145832 423678 145888
rect 423734 145832 423739 145888
rect 377949 145830 423739 145832
rect 377949 145827 378015 145830
rect 423673 145827 423739 145830
rect 56317 145754 56383 145757
rect 99373 145754 99439 145757
rect 56317 145752 99439 145754
rect 56317 145696 56322 145752
rect 56378 145696 99378 145752
rect 99434 145696 99439 145752
rect 56317 145694 99439 145696
rect 56317 145691 56383 145694
rect 99373 145691 99439 145694
rect 370313 145754 370379 145757
rect 377806 145754 377812 145756
rect 370313 145752 377812 145754
rect 370313 145696 370318 145752
rect 370374 145696 377812 145752
rect 370313 145694 377812 145696
rect 370313 145691 370379 145694
rect 377806 145692 377812 145694
rect 377876 145754 377882 145756
rect 425053 145754 425119 145757
rect 377876 145752 425119 145754
rect 377876 145696 425058 145752
rect 425114 145696 425119 145752
rect 377876 145694 425119 145696
rect 377876 145692 377882 145694
rect 425053 145691 425119 145694
rect 50245 145618 50311 145621
rect 54569 145618 54635 145621
rect 98637 145618 98703 145621
rect 50245 145616 98703 145618
rect 50245 145560 50250 145616
rect 50306 145560 54574 145616
rect 54630 145560 98642 145616
rect 98698 145560 98703 145616
rect 50245 145558 98703 145560
rect 50245 145555 50311 145558
rect 54569 145555 54635 145558
rect 98637 145555 98703 145558
rect 213453 145618 213519 145621
rect 237373 145618 237439 145621
rect 213453 145616 237439 145618
rect 213453 145560 213458 145616
rect 213514 145560 237378 145616
rect 237434 145560 237439 145616
rect 213453 145558 237439 145560
rect 213453 145555 213519 145558
rect 237373 145555 237439 145558
rect 369761 145618 369827 145621
rect 377489 145618 377555 145621
rect 377949 145618 378015 145621
rect 369761 145616 378015 145618
rect 369761 145560 369766 145616
rect 369822 145560 377494 145616
rect 377550 145560 377954 145616
rect 378010 145560 378015 145616
rect 369761 145558 378015 145560
rect 369761 145555 369827 145558
rect 377489 145555 377555 145558
rect 377949 145555 378015 145558
rect 379462 145556 379468 145620
rect 379532 145618 379538 145620
rect 429193 145618 429259 145621
rect 379532 145616 429259 145618
rect 379532 145560 429198 145616
rect 429254 145560 429259 145616
rect 379532 145558 429259 145560
rect 379532 145556 379538 145558
rect 429193 145555 429259 145558
rect 510613 145482 510679 145485
rect 510838 145482 510844 145484
rect 510613 145480 510844 145482
rect 510613 145424 510618 145480
rect 510674 145424 510844 145480
rect 510613 145422 510844 145424
rect 510613 145419 510679 145422
rect 510838 145420 510844 145422
rect 510908 145420 510914 145484
rect 178534 144876 178540 144940
rect 178604 144938 178610 144940
rect 179045 144938 179111 144941
rect 179689 144940 179755 144941
rect 179638 144938 179644 144940
rect 178604 144936 179111 144938
rect 178604 144880 179050 144936
rect 179106 144880 179111 144936
rect 178604 144878 179111 144880
rect 179598 144878 179644 144938
rect 179708 144936 179755 144940
rect 179750 144880 179755 144936
rect 178604 144876 178610 144878
rect 179045 144875 179111 144878
rect 179638 144876 179644 144878
rect 179708 144876 179755 144880
rect 190862 144876 190868 144940
rect 190932 144938 190938 144940
rect 191281 144938 191347 144941
rect 338481 144940 338547 144941
rect 338430 144938 338436 144940
rect 190932 144936 191347 144938
rect 190932 144880 191286 144936
rect 191342 144880 191347 144936
rect 190932 144878 191347 144880
rect 338390 144878 338436 144938
rect 338500 144936 338547 144940
rect 338542 144880 338547 144936
rect 190932 144876 190938 144878
rect 179689 144875 179755 144876
rect 191281 144875 191347 144878
rect 338430 144876 338436 144878
rect 338500 144876 338547 144880
rect 339718 144876 339724 144940
rect 339788 144938 339794 144940
rect 340229 144938 340295 144941
rect 339788 144936 340295 144938
rect 339788 144880 340234 144936
rect 340290 144880 340295 144936
rect 339788 144878 340295 144880
rect 339788 144876 339794 144878
rect 338481 144875 338547 144876
rect 340229 144875 340295 144878
rect 350942 144876 350948 144940
rect 351012 144938 351018 144940
rect 351637 144938 351703 144941
rect 351012 144936 351703 144938
rect 351012 144880 351642 144936
rect 351698 144880 351703 144936
rect 351012 144878 351703 144880
rect 351012 144876 351018 144878
rect 351637 144875 351703 144878
rect 498510 144876 498516 144940
rect 498580 144938 498586 144940
rect 498653 144938 498719 144941
rect 498580 144936 498719 144938
rect 498580 144880 498658 144936
rect 498714 144880 498719 144936
rect 498580 144878 498719 144880
rect 498580 144876 498586 144878
rect 498653 144875 498719 144878
rect 499798 144876 499804 144940
rect 499868 144938 499874 144940
rect 500217 144938 500283 144941
rect 499868 144936 500283 144938
rect 499868 144880 500222 144936
rect 500278 144880 500283 144936
rect 499868 144878 500283 144880
rect 499868 144876 499874 144878
rect 500217 144875 500283 144878
rect 57462 140796 57468 140860
rect 57532 140858 57538 140860
rect 59445 140858 59511 140861
rect 57532 140856 59511 140858
rect 57532 140800 59450 140856
rect 59506 140800 59511 140856
rect 57532 140798 59511 140800
rect 57532 140796 57538 140798
rect 59445 140795 59511 140798
rect 358905 139362 358971 139365
rect 519077 139362 519143 139365
rect 356562 139360 358971 139362
rect 356562 139304 358910 139360
rect 358966 139304 358971 139360
rect 356562 139302 358971 139304
rect 198825 139226 198891 139229
rect 197126 139224 198891 139226
rect 197126 139220 198830 139224
rect 196604 139168 198830 139220
rect 198886 139168 198891 139224
rect 356562 139190 356622 139302
rect 358905 139299 358971 139302
rect 516558 139360 519143 139362
rect 516558 139304 519082 139360
rect 519138 139304 519143 139360
rect 516558 139302 519143 139304
rect 516558 139190 516618 139302
rect 519077 139299 519143 139302
rect 583520 139212 584960 139452
rect 196604 139166 198891 139168
rect 196604 139160 197186 139166
rect 198825 139163 198891 139166
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 57145 97474 57211 97477
rect 57145 97472 60062 97474
rect 57145 97416 57150 97472
rect 57206 97416 60062 97472
rect 57145 97414 60062 97416
rect 57145 97411 57211 97414
rect 60002 96894 60062 97414
rect 217409 96930 217475 96933
rect 377305 96930 377371 96933
rect 217409 96928 219450 96930
rect 217409 96872 217414 96928
rect 217470 96924 219450 96928
rect 377305 96928 379530 96930
rect 217470 96872 220064 96924
rect 217409 96870 220064 96872
rect 217409 96867 217475 96870
rect 219390 96864 220064 96870
rect 377305 96872 377310 96928
rect 377366 96924 379530 96928
rect 377366 96872 380052 96924
rect 377305 96870 380052 96872
rect 377305 96867 377371 96870
rect 379470 96864 380052 96870
rect 56777 96522 56843 96525
rect 56777 96520 60062 96522
rect 56777 96464 56782 96520
rect 56838 96464 60062 96520
rect 56777 96462 60062 96464
rect 56777 96459 56843 96462
rect 60002 95942 60062 96462
rect 217593 95978 217659 95981
rect 377029 95978 377095 95981
rect 217593 95976 219450 95978
rect 217593 95920 217598 95976
rect 217654 95972 219450 95976
rect 377029 95976 379530 95978
rect 217654 95920 220064 95972
rect 217593 95918 220064 95920
rect 217593 95915 217659 95918
rect 219390 95912 220064 95918
rect 377029 95920 377034 95976
rect 377090 95972 379530 95976
rect 377090 95920 380052 95972
rect 377029 95918 380052 95920
rect 377029 95915 377095 95918
rect 379470 95912 380052 95918
rect 57605 93802 57671 93805
rect 217685 93802 217751 93805
rect 376937 93802 377003 93805
rect 57605 93800 60062 93802
rect 57605 93744 57610 93800
rect 57666 93744 60062 93800
rect 57605 93742 60062 93744
rect 217685 93800 219450 93802
rect 217685 93744 217690 93800
rect 217746 93796 219450 93800
rect 376937 93800 379530 93802
rect 217746 93744 220064 93796
rect 217685 93742 220064 93744
rect 57605 93739 57671 93742
rect 217685 93739 217751 93742
rect 219390 93736 220064 93742
rect 376937 93744 376942 93800
rect 376998 93796 379530 93800
rect 376998 93744 380052 93796
rect 376937 93742 380052 93744
rect 376937 93739 377003 93742
rect 379470 93736 380052 93742
rect 57329 93394 57395 93397
rect 57329 93392 60062 93394
rect 57329 93336 57334 93392
rect 57390 93336 60062 93392
rect 57329 93334 60062 93336
rect 57329 93331 57395 93334
rect 60002 92814 60062 93334
rect 217225 92850 217291 92853
rect 377213 92850 377279 92853
rect 217225 92848 219450 92850
rect 217225 92792 217230 92848
rect 217286 92844 219450 92848
rect 377213 92848 379530 92850
rect 217286 92792 220064 92844
rect 217225 92790 220064 92792
rect 217225 92787 217291 92790
rect 219390 92784 220064 92790
rect 377213 92792 377218 92848
rect 377274 92844 379530 92848
rect 377274 92792 380052 92844
rect 377213 92790 380052 92792
rect 377213 92787 377279 92790
rect 379470 92784 380052 92790
rect 57789 91082 57855 91085
rect 217501 91082 217567 91085
rect 377673 91082 377739 91085
rect 57789 91080 60062 91082
rect 57789 91024 57794 91080
rect 57850 91024 60062 91080
rect 57789 91022 60062 91024
rect 217501 91080 219450 91082
rect 217501 91024 217506 91080
rect 217562 91076 219450 91080
rect 377673 91080 379530 91082
rect 217562 91024 220064 91076
rect 217501 91022 220064 91024
rect 57789 91019 57855 91022
rect 217501 91019 217567 91022
rect 219390 91016 220064 91022
rect 377673 91024 377678 91080
rect 377734 91076 379530 91080
rect 377734 91024 380052 91076
rect 377673 91022 380052 91024
rect 377673 91019 377739 91022
rect 379470 91016 380052 91022
rect 57421 90538 57487 90541
rect 57421 90536 60062 90538
rect 57421 90480 57426 90536
rect 57482 90480 60062 90536
rect 57421 90478 60062 90480
rect 57421 90475 57487 90478
rect 60002 89958 60062 90478
rect 216765 89994 216831 89997
rect 377857 89994 377923 89997
rect 216765 89992 219450 89994
rect 216765 89936 216770 89992
rect 216826 89988 219450 89992
rect 377857 89992 379530 89994
rect 216826 89936 220064 89988
rect 216765 89934 220064 89936
rect 216765 89931 216831 89934
rect 219390 89928 220064 89934
rect 377857 89936 377862 89992
rect 377918 89988 379530 89992
rect 377918 89936 380052 89988
rect 377857 89934 380052 89936
rect 377857 89931 377923 89934
rect 379470 89928 380052 89934
rect 57697 88226 57763 88229
rect 217777 88226 217843 88229
rect 377765 88226 377831 88229
rect 57697 88224 60062 88226
rect 57697 88168 57702 88224
rect 57758 88168 60062 88224
rect 57697 88166 60062 88168
rect 217777 88224 219450 88226
rect 217777 88168 217782 88224
rect 217838 88220 219450 88224
rect 377765 88224 379530 88226
rect 217838 88168 220064 88220
rect 217777 88166 220064 88168
rect 57697 88163 57763 88166
rect 217777 88163 217843 88166
rect 219390 88160 220064 88166
rect 377765 88168 377770 88224
rect 377826 88220 379530 88224
rect 377826 88168 380052 88220
rect 377765 88166 380052 88168
rect 377765 88163 377831 88166
rect 379470 88160 380052 88166
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 359457 79930 359523 79933
rect 518893 79930 518959 79933
rect 520181 79930 520247 79933
rect 356562 79928 359523 79930
rect 356562 79872 359462 79928
rect 359518 79872 359523 79928
rect 356562 79870 359523 79872
rect 199285 79386 199351 79389
rect 197126 79384 199351 79386
rect 197126 79380 199290 79384
rect 196604 79328 199290 79380
rect 199346 79328 199351 79384
rect 356562 79350 356622 79870
rect 359457 79867 359523 79870
rect 516558 79928 520247 79930
rect 516558 79872 518898 79928
rect 518954 79872 520186 79928
rect 520242 79872 520247 79928
rect 516558 79870 520247 79872
rect 516558 79350 516618 79870
rect 518893 79867 518959 79870
rect 520181 79867 520247 79870
rect 196604 79326 199351 79328
rect 196604 79320 197186 79326
rect 199285 79323 199351 79326
rect 359365 78298 359431 78301
rect 519445 78298 519511 78301
rect 356562 78296 359431 78298
rect 356562 78240 359370 78296
rect 359426 78240 359431 78296
rect 356562 78238 359431 78240
rect 199193 77754 199259 77757
rect 197126 77752 199259 77754
rect 197126 77748 199198 77752
rect 196604 77696 199198 77748
rect 199254 77696 199259 77752
rect 356562 77718 356622 78238
rect 359365 78235 359431 78238
rect 516558 78296 519511 78298
rect 516558 78240 519450 78296
rect 519506 78240 519511 78296
rect 516558 78238 519511 78240
rect 516558 77718 516618 78238
rect 519445 78235 519511 78238
rect 196604 77694 199259 77696
rect 196604 77688 197186 77694
rect 199193 77691 199259 77694
rect 359181 76938 359247 76941
rect 356562 76936 359247 76938
rect 356562 76880 359186 76936
rect 359242 76880 359247 76936
rect 356562 76878 359247 76880
rect 198917 76394 198983 76397
rect 197126 76392 198983 76394
rect 197126 76388 198922 76392
rect 196604 76336 198922 76388
rect 198978 76336 198983 76392
rect 356562 76358 356622 76878
rect 359181 76875 359247 76878
rect 519353 76802 519419 76805
rect 516558 76800 519419 76802
rect 516558 76744 519358 76800
rect 519414 76744 519419 76800
rect 516558 76742 519419 76744
rect 516558 76358 516618 76742
rect 519353 76739 519419 76742
rect 196604 76334 198983 76336
rect 196604 76328 197186 76334
rect 198917 76331 198983 76334
rect 359089 75442 359155 75445
rect 518985 75442 519051 75445
rect 356562 75440 359155 75442
rect 356562 75384 359094 75440
rect 359150 75384 359155 75440
rect 356562 75382 359155 75384
rect 198733 74898 198799 74901
rect 197126 74896 198799 74898
rect 197126 74892 198738 74896
rect 196604 74840 198738 74892
rect 198794 74840 198799 74896
rect 356562 74862 356622 75382
rect 359089 75379 359155 75382
rect 516558 75440 519051 75442
rect 516558 75384 518990 75440
rect 519046 75384 519051 75440
rect 516558 75382 519051 75384
rect 516558 74862 516618 75382
rect 518985 75379 519051 75382
rect 196604 74838 198799 74840
rect 196604 74832 197186 74838
rect 198733 74835 198799 74838
rect 519169 74218 519235 74221
rect 516558 74216 519235 74218
rect 516558 74160 519174 74216
rect 519230 74160 519235 74216
rect 516558 74158 519235 74160
rect 359273 74082 359339 74085
rect 356562 74080 359339 74082
rect 356562 74024 359278 74080
rect 359334 74024 359339 74080
rect 356562 74022 359339 74024
rect 199009 73674 199075 73677
rect 197126 73672 199075 73674
rect 197126 73668 199014 73672
rect 196604 73616 199014 73668
rect 199070 73616 199075 73672
rect 356562 73638 356622 74022
rect 359273 74019 359339 74022
rect 516558 73638 516618 74158
rect 519169 74155 519235 74158
rect 196604 73614 199075 73616
rect 196604 73608 197186 73614
rect 199009 73611 199075 73614
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 57605 70138 57671 70141
rect 57605 70136 60062 70138
rect 57605 70080 57610 70136
rect 57666 70080 60062 70136
rect 57605 70078 60062 70080
rect 57605 70075 57671 70078
rect 60002 69966 60062 70078
rect 216673 70002 216739 70005
rect 376937 70002 377003 70005
rect 216673 70000 219450 70002
rect 216673 69944 216678 70000
rect 216734 69996 219450 70000
rect 376937 70000 379530 70002
rect 216734 69944 220064 69996
rect 216673 69942 220064 69944
rect 216673 69939 216739 69942
rect 219390 69936 220064 69942
rect 376937 69944 376942 70000
rect 376998 69996 379530 70000
rect 376998 69944 380052 69996
rect 376937 69942 380052 69944
rect 376937 69939 377003 69942
rect 379470 69936 380052 69942
rect 57881 68914 57947 68917
rect 57881 68912 60062 68914
rect 57881 68856 57886 68912
rect 57942 68856 60062 68912
rect 57881 68854 60062 68856
rect 57881 68851 57947 68854
rect 60002 68334 60062 68854
rect 216673 68370 216739 68373
rect 217961 68370 218027 68373
rect 376937 68370 377003 68373
rect 216673 68368 219450 68370
rect 216673 68312 216678 68368
rect 216734 68312 217966 68368
rect 218022 68364 219450 68368
rect 376937 68368 379530 68370
rect 218022 68312 220064 68364
rect 216673 68310 220064 68312
rect 216673 68307 216739 68310
rect 217961 68307 218027 68310
rect 219390 68304 220064 68310
rect 376937 68312 376942 68368
rect 376998 68364 379530 68368
rect 376998 68312 380052 68364
rect 376937 68310 380052 68312
rect 376937 68307 377003 68310
rect 379470 68304 380052 68310
rect 46790 67764 46796 67828
rect 46860 67826 46866 67828
rect 60002 67826 60062 68062
rect 214414 68036 214420 68100
rect 214484 68098 214490 68100
rect 214484 68092 219450 68098
rect 214484 68038 220064 68092
rect 214484 68036 214490 68038
rect 219390 68032 220064 68038
rect 376150 68036 376156 68100
rect 376220 68098 376226 68100
rect 376220 68092 379530 68098
rect 376220 68038 380052 68092
rect 376220 68036 376226 68038
rect 379470 68032 380052 68038
rect 46860 67766 60062 67826
rect 46860 67764 46866 67766
rect 219065 60620 219131 60621
rect 219014 60618 219020 60620
rect 218974 60558 219020 60618
rect 219084 60616 219131 60620
rect 219126 60560 219131 60616
rect 219014 60556 219020 60558
rect 219084 60556 219131 60560
rect 219065 60555 219131 60556
rect 77109 59804 77175 59805
rect 83089 59804 83155 59805
rect 101765 59804 101831 59805
rect 77109 59800 77142 59804
rect 77206 59802 77212 59804
rect 77109 59744 77114 59800
rect 77109 59740 77142 59744
rect 77206 59742 77266 59802
rect 83089 59800 83126 59804
rect 83190 59802 83196 59804
rect 101752 59802 101758 59804
rect 83089 59744 83094 59800
rect 77206 59740 77212 59742
rect 83089 59740 83126 59744
rect 83190 59742 83246 59802
rect 101674 59742 101758 59802
rect 101822 59800 101831 59804
rect 101826 59744 101831 59800
rect 83190 59740 83196 59742
rect 101752 59740 101758 59742
rect 101822 59740 101831 59744
rect 77109 59739 77175 59740
rect 83089 59739 83155 59740
rect 101765 59739 101831 59740
rect 103881 59804 103947 59805
rect 107561 59804 107627 59805
rect 113541 59804 113607 59805
rect 235993 59804 236059 59805
rect 237097 59804 237163 59805
rect 255865 59804 255931 59805
rect 256969 59804 257035 59805
rect 262857 59804 262923 59805
rect 396073 59804 396139 59805
rect 103881 59800 103934 59804
rect 103998 59802 104004 59804
rect 103881 59744 103886 59800
rect 103881 59740 103934 59744
rect 103998 59742 104038 59802
rect 107561 59800 107606 59804
rect 107670 59802 107676 59804
rect 107561 59744 107566 59800
rect 103998 59740 104004 59742
rect 107561 59740 107606 59744
rect 107670 59742 107718 59802
rect 113541 59800 113590 59804
rect 113654 59802 113660 59804
rect 113541 59744 113546 59800
rect 107670 59740 107676 59742
rect 113541 59740 113590 59744
rect 113654 59742 113698 59802
rect 235993 59800 236054 59804
rect 235993 59744 235998 59800
rect 113654 59740 113660 59742
rect 235993 59740 236054 59744
rect 236118 59802 236124 59804
rect 236118 59742 236150 59802
rect 237097 59800 237142 59804
rect 237206 59802 237212 59804
rect 237097 59744 237102 59800
rect 236118 59740 236124 59742
rect 237097 59740 237142 59744
rect 237206 59742 237254 59802
rect 255865 59800 255910 59804
rect 255974 59802 255980 59804
rect 255865 59744 255870 59800
rect 237206 59740 237212 59742
rect 255865 59740 255910 59744
rect 255974 59742 256022 59802
rect 256969 59800 256998 59804
rect 257062 59802 257068 59804
rect 262840 59802 262846 59804
rect 256969 59744 256974 59800
rect 255974 59740 255980 59742
rect 256969 59740 256998 59744
rect 257062 59742 257126 59802
rect 262766 59742 262846 59802
rect 262910 59800 262923 59804
rect 396048 59802 396054 59804
rect 262918 59744 262923 59800
rect 257062 59740 257068 59742
rect 262840 59740 262846 59742
rect 262910 59740 262923 59744
rect 395982 59742 396054 59802
rect 396118 59800 396139 59804
rect 396134 59744 396139 59800
rect 396048 59740 396054 59742
rect 396118 59740 396139 59744
rect 103881 59739 103947 59740
rect 107561 59739 107627 59740
rect 113541 59739 113607 59740
rect 235993 59739 236059 59740
rect 237097 59739 237163 59740
rect 255865 59739 255931 59740
rect 256969 59739 257035 59740
rect 262857 59739 262923 59740
rect 396073 59739 396139 59740
rect 397085 59804 397151 59805
rect 403065 59804 403131 59805
rect 416957 59804 417023 59805
rect 422845 59804 422911 59805
rect 423949 59804 424015 59805
rect 397085 59800 397142 59804
rect 397206 59802 397212 59804
rect 397085 59744 397090 59800
rect 397085 59740 397142 59744
rect 397206 59742 397242 59802
rect 403065 59800 403126 59804
rect 403065 59744 403070 59800
rect 397206 59740 397212 59742
rect 403065 59740 403126 59744
rect 403190 59802 403196 59804
rect 403190 59742 403222 59802
rect 416957 59800 416998 59804
rect 417062 59802 417068 59804
rect 422840 59802 422846 59804
rect 416957 59744 416962 59800
rect 403190 59740 403196 59742
rect 416957 59740 416998 59744
rect 417062 59742 417114 59802
rect 422754 59742 422846 59802
rect 417062 59740 417068 59742
rect 422840 59740 422846 59742
rect 422910 59740 422916 59804
rect 423928 59802 423934 59804
rect 423858 59742 423934 59802
rect 423998 59800 424015 59804
rect 424010 59744 424015 59800
rect 423928 59740 423934 59742
rect 423998 59740 424015 59744
rect 397085 59739 397151 59740
rect 403065 59739 403131 59740
rect 416957 59739 417023 59740
rect 422845 59739 422911 59740
rect 423949 59739 424015 59740
rect 94497 59668 94563 59669
rect 96981 59668 97047 59669
rect 98085 59668 98151 59669
rect 100753 59668 100819 59669
rect 94497 59664 94550 59668
rect 94614 59666 94620 59668
rect 94497 59608 94502 59664
rect 94497 59604 94550 59608
rect 94614 59606 94654 59666
rect 96981 59664 96998 59668
rect 97062 59666 97068 59668
rect 98080 59666 98086 59668
rect 96981 59608 96986 59664
rect 94614 59604 94620 59606
rect 96981 59604 96998 59608
rect 97062 59606 97138 59666
rect 97994 59606 98086 59666
rect 97062 59604 97068 59606
rect 98080 59604 98086 59606
rect 98150 59604 98156 59668
rect 100702 59666 100708 59668
rect 100662 59606 100708 59666
rect 100772 59664 100819 59668
rect 100814 59608 100819 59664
rect 100702 59604 100708 59606
rect 100772 59604 100819 59608
rect 94497 59603 94563 59604
rect 96981 59603 97047 59604
rect 98085 59603 98151 59604
rect 100753 59603 100819 59604
rect 102777 59668 102843 59669
rect 108665 59668 108731 59669
rect 260649 59668 260715 59669
rect 308489 59668 308555 59669
rect 315849 59668 315915 59669
rect 404169 59668 404235 59669
rect 102777 59664 102846 59668
rect 102777 59608 102782 59664
rect 102838 59608 102846 59664
rect 102777 59604 102846 59608
rect 102910 59666 102916 59668
rect 105968 59666 105974 59668
rect 102910 59606 102934 59666
rect 103470 59606 105974 59666
rect 102910 59604 102916 59606
rect 102777 59603 102843 59604
rect 95877 59532 95943 59533
rect 95877 59528 95924 59532
rect 95988 59530 95994 59532
rect 95877 59472 95882 59528
rect 95877 59468 95924 59472
rect 95988 59470 96034 59530
rect 95988 59468 95994 59470
rect 95877 59467 95943 59468
rect 46606 59332 46612 59396
rect 46676 59394 46682 59396
rect 103470 59394 103530 59606
rect 105968 59604 105974 59606
rect 106038 59604 106044 59668
rect 108665 59664 108694 59668
rect 108758 59666 108764 59668
rect 108665 59608 108670 59664
rect 108665 59604 108694 59608
rect 108758 59606 108822 59666
rect 260649 59664 260670 59668
rect 260734 59666 260740 59668
rect 260649 59608 260654 59664
rect 108758 59604 108764 59606
rect 260649 59604 260670 59608
rect 260734 59606 260806 59666
rect 308489 59664 308542 59668
rect 308606 59666 308612 59668
rect 308489 59608 308494 59664
rect 260734 59604 260740 59606
rect 308489 59604 308542 59608
rect 308606 59606 308646 59666
rect 315849 59664 315886 59668
rect 315950 59666 315956 59668
rect 315849 59608 315854 59664
rect 308606 59604 308612 59606
rect 315849 59604 315886 59608
rect 315950 59606 316006 59666
rect 404169 59664 404214 59668
rect 404278 59666 404284 59668
rect 412541 59666 412607 59669
rect 423489 59668 423555 59669
rect 413456 59666 413462 59668
rect 404169 59608 404174 59664
rect 315950 59604 315956 59606
rect 404169 59604 404214 59608
rect 404278 59606 404326 59666
rect 412541 59664 413462 59666
rect 412541 59608 412546 59664
rect 412602 59608 413462 59664
rect 412541 59606 413462 59608
rect 404278 59604 404284 59606
rect 108665 59603 108731 59604
rect 260649 59603 260715 59604
rect 308489 59603 308555 59604
rect 315849 59603 315915 59604
rect 404169 59603 404235 59604
rect 412541 59603 412607 59606
rect 413456 59604 413462 59606
rect 413526 59604 413532 59668
rect 423489 59664 423526 59668
rect 423590 59666 423596 59668
rect 423489 59608 423494 59664
rect 423489 59604 423526 59608
rect 423590 59606 423646 59666
rect 423590 59604 423596 59606
rect 423489 59603 423555 59604
rect 263542 59530 263548 59532
rect 258030 59470 263548 59530
rect 46676 59334 103530 59394
rect 110965 59396 111031 59397
rect 110965 59392 111012 59396
rect 111076 59394 111082 59396
rect 110965 59336 110970 59392
rect 46676 59332 46682 59334
rect 110965 59332 111012 59336
rect 111076 59334 111122 59394
rect 111076 59332 111082 59334
rect 200798 59332 200804 59396
rect 200868 59394 200874 59396
rect 258030 59394 258090 59470
rect 263542 59468 263548 59470
rect 263612 59468 263618 59532
rect 583520 59516 584960 59756
rect 200868 59334 258090 59394
rect 259453 59396 259519 59397
rect 261661 59396 261727 59397
rect 410701 59396 410767 59397
rect 414565 59396 414631 59397
rect 416037 59396 416103 59397
rect 418153 59396 418219 59397
rect 259453 59392 259500 59396
rect 259564 59394 259570 59396
rect 259453 59336 259458 59392
rect 200868 59332 200874 59334
rect 259453 59332 259500 59336
rect 259564 59334 259610 59394
rect 261661 59392 261708 59396
rect 261772 59394 261778 59396
rect 261661 59336 261666 59392
rect 259564 59332 259570 59334
rect 261661 59332 261708 59336
rect 261772 59334 261818 59394
rect 410701 59392 410748 59396
rect 410812 59394 410818 59396
rect 410701 59336 410706 59392
rect 261772 59332 261778 59334
rect 410701 59332 410748 59336
rect 410812 59334 410858 59394
rect 414565 59392 414612 59396
rect 414676 59394 414682 59396
rect 414565 59336 414570 59392
rect 410812 59332 410818 59334
rect 414565 59332 414612 59336
rect 414676 59334 414722 59394
rect 416037 59392 416084 59396
rect 416148 59394 416154 59396
rect 418102 59394 418108 59396
rect 416037 59336 416042 59392
rect 414676 59332 414682 59334
rect 416037 59332 416084 59336
rect 416148 59334 416194 59394
rect 418062 59334 418108 59394
rect 418172 59392 418219 59396
rect 418214 59336 418219 59392
rect 416148 59332 416154 59334
rect 418102 59332 418108 59334
rect 418172 59332 418219 59336
rect 110965 59331 111031 59332
rect 259453 59331 259519 59332
rect 261661 59331 261727 59332
rect 410701 59331 410767 59332
rect 414565 59331 414631 59332
rect 416037 59331 416103 59332
rect 418153 59331 418219 59332
rect 419349 59396 419415 59397
rect 420637 59396 420703 59397
rect 421741 59396 421807 59397
rect 428181 59396 428247 59397
rect 419349 59392 419396 59396
rect 419460 59394 419466 59396
rect 419349 59336 419354 59392
rect 419349 59332 419396 59336
rect 419460 59334 419506 59394
rect 420637 59392 420684 59396
rect 420748 59394 420754 59396
rect 420637 59336 420642 59392
rect 419460 59332 419466 59334
rect 420637 59332 420684 59336
rect 420748 59334 420794 59394
rect 421741 59392 421788 59396
rect 421852 59394 421858 59396
rect 421741 59336 421746 59392
rect 420748 59332 420754 59334
rect 421741 59332 421788 59336
rect 421852 59334 421898 59394
rect 428181 59392 428228 59396
rect 428292 59394 428298 59396
rect 428181 59336 428186 59392
rect 421852 59332 421858 59334
rect 428181 59332 428228 59336
rect 428292 59334 428338 59394
rect 428292 59332 428298 59334
rect 419349 59331 419415 59332
rect 420637 59331 420703 59332
rect 421741 59331 421807 59332
rect 428181 59331 428247 59332
rect 148501 59260 148567 59261
rect 150893 59260 150959 59261
rect 279233 59260 279299 59261
rect 54886 59196 54892 59260
rect 54956 59258 54962 59260
rect 143574 59258 143580 59260
rect 54956 59198 143580 59258
rect 54956 59196 54962 59198
rect 143574 59196 143580 59198
rect 143644 59196 143650 59260
rect 148501 59256 148548 59260
rect 148612 59258 148618 59260
rect 148501 59200 148506 59256
rect 148501 59196 148548 59200
rect 148612 59198 148658 59258
rect 150893 59256 150940 59260
rect 151004 59258 151010 59260
rect 150893 59200 150898 59256
rect 148612 59196 148618 59198
rect 150893 59196 150940 59200
rect 151004 59198 151050 59258
rect 151004 59196 151010 59198
rect 198406 59196 198412 59260
rect 198476 59258 198482 59260
rect 276054 59258 276060 59260
rect 198476 59198 276060 59258
rect 198476 59196 198482 59198
rect 276054 59196 276060 59198
rect 276124 59196 276130 59260
rect 279182 59258 279188 59260
rect 279142 59198 279188 59258
rect 279252 59256 279299 59260
rect 279294 59200 279299 59256
rect 279182 59196 279188 59198
rect 279252 59196 279299 59200
rect 148501 59195 148567 59196
rect 150893 59195 150959 59196
rect 279233 59195 279299 59196
rect 290917 59260 290983 59261
rect 300853 59260 300919 59261
rect 320909 59260 320975 59261
rect 325877 59260 325943 59261
rect 290917 59256 290964 59260
rect 291028 59258 291034 59260
rect 290917 59200 290922 59256
rect 290917 59196 290964 59200
rect 291028 59198 291074 59258
rect 300853 59256 300900 59260
rect 300964 59258 300970 59260
rect 300853 59200 300858 59256
rect 291028 59196 291034 59198
rect 300853 59196 300900 59200
rect 300964 59198 301010 59258
rect 320909 59256 320956 59260
rect 321020 59258 321026 59260
rect 320909 59200 320914 59256
rect 300964 59196 300970 59198
rect 320909 59196 320956 59200
rect 321020 59198 321066 59258
rect 325877 59256 325924 59260
rect 325988 59258 325994 59260
rect 325877 59200 325882 59256
rect 321020 59196 321026 59198
rect 325877 59196 325924 59200
rect 325988 59198 326034 59258
rect 325988 59196 325994 59198
rect 357934 59196 357940 59260
rect 358004 59258 358010 59260
rect 480846 59258 480852 59260
rect 358004 59198 480852 59258
rect 358004 59196 358010 59198
rect 480846 59196 480852 59198
rect 480916 59196 480922 59260
rect 290917 59195 290983 59196
rect 300853 59195 300919 59196
rect 320909 59195 320975 59196
rect 325877 59195 325943 59196
rect 53414 59060 53420 59124
rect 53484 59122 53490 59124
rect 140814 59122 140820 59124
rect 53484 59062 140820 59122
rect 53484 59060 53490 59062
rect 140814 59060 140820 59062
rect 140884 59060 140890 59124
rect 206870 59060 206876 59124
rect 206940 59122 206946 59124
rect 280838 59122 280844 59124
rect 206940 59062 280844 59122
rect 206940 59060 206946 59062
rect 280838 59060 280844 59062
rect 280908 59060 280914 59124
rect 373758 59060 373764 59124
rect 373828 59122 373834 59124
rect 483422 59122 483428 59124
rect 373828 59062 483428 59122
rect 373828 59060 373834 59062
rect 483422 59060 483428 59062
rect 483492 59060 483498 59124
rect 475837 58988 475903 58989
rect 52126 58924 52132 58988
rect 52196 58986 52202 58988
rect 138422 58986 138428 58988
rect 52196 58926 138428 58986
rect 52196 58924 52202 58926
rect 138422 58924 138428 58926
rect 138492 58924 138498 58988
rect 212390 58924 212396 58988
rect 212460 58986 212466 58988
rect 285990 58986 285996 58988
rect 212460 58926 285996 58986
rect 212460 58924 212466 58926
rect 285990 58924 285996 58926
rect 286060 58924 286066 58988
rect 371734 58924 371740 58988
rect 371804 58986 371810 58988
rect 473486 58986 473492 58988
rect 371804 58926 473492 58986
rect 371804 58924 371810 58926
rect 473486 58924 473492 58926
rect 473556 58924 473562 58988
rect 475837 58984 475884 58988
rect 475948 58986 475954 58988
rect 475837 58928 475842 58984
rect 475837 58924 475884 58928
rect 475948 58926 475994 58986
rect 475948 58924 475954 58926
rect 475837 58923 475903 58924
rect 468477 58852 468543 58853
rect 55438 58788 55444 58852
rect 55508 58850 55514 58852
rect 135846 58850 135852 58852
rect 55508 58790 135852 58850
rect 55508 58788 55514 58790
rect 135846 58788 135852 58790
rect 135916 58788 135922 58852
rect 198590 58788 198596 58852
rect 198660 58850 198666 58852
rect 268326 58850 268332 58852
rect 198660 58790 268332 58850
rect 198660 58788 198666 58790
rect 268326 58788 268332 58790
rect 268396 58788 268402 58852
rect 364926 58788 364932 58852
rect 364996 58850 365002 58852
rect 453430 58850 453436 58852
rect 364996 58790 453436 58850
rect 364996 58788 365002 58790
rect 453430 58788 453436 58790
rect 453500 58788 453506 58852
rect 468477 58848 468524 58852
rect 468588 58850 468594 58852
rect 468477 58792 468482 58848
rect 468477 58788 468524 58792
rect 468588 58790 468634 58850
rect 468588 58788 468594 58790
rect 468477 58787 468543 58788
rect -960 58578 480 58668
rect 59302 58652 59308 58716
rect 59372 58714 59378 58716
rect 120942 58714 120948 58716
rect 59372 58654 120948 58714
rect 59372 58652 59378 58654
rect 120942 58652 120948 58654
rect 121012 58652 121018 58716
rect 197854 58652 197860 58716
rect 197924 58714 197930 58716
rect 253606 58714 253612 58716
rect 197924 58654 253612 58714
rect 197924 58652 197930 58654
rect 253606 58652 253612 58654
rect 253676 58652 253682 58716
rect 374494 58652 374500 58716
rect 374564 58714 374570 58716
rect 463550 58714 463556 58716
rect 374564 58654 463556 58714
rect 374564 58652 374570 58654
rect 463550 58652 463556 58654
rect 463620 58652 463626 58716
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 48078 58516 48084 58580
rect 48148 58578 48154 58580
rect 108246 58578 108252 58580
rect 48148 58518 108252 58578
rect 48148 58516 48154 58518
rect 108246 58516 108252 58518
rect 108316 58516 108322 58580
rect 200614 58516 200620 58580
rect 200684 58578 200690 58580
rect 250662 58578 250668 58580
rect 200684 58518 250668 58578
rect 200684 58516 200690 58518
rect 250662 58516 250668 58518
rect 250732 58516 250738 58580
rect 375966 58516 375972 58580
rect 376036 58578 376042 58580
rect 458398 58578 458404 58580
rect 376036 58518 458404 58578
rect 376036 58516 376042 58518
rect 458398 58516 458404 58518
rect 458468 58516 458474 58580
rect 59118 58380 59124 58444
rect 59188 58442 59194 58444
rect 101070 58442 101076 58444
rect 59188 58382 101076 58442
rect 59188 58380 59194 58382
rect 101070 58380 101076 58382
rect 101140 58380 101146 58444
rect 217542 58380 217548 58444
rect 217612 58442 217618 58444
rect 257838 58442 257844 58444
rect 217612 58382 257844 58442
rect 217612 58380 217618 58382
rect 257838 58380 257844 58382
rect 257908 58380 257914 58444
rect 85430 58108 85436 58172
rect 85500 58108 85506 58172
rect 92238 58108 92244 58172
rect 92308 58108 92314 58172
rect 99414 58108 99420 58172
rect 99484 58108 99490 58172
rect 128302 58108 128308 58172
rect 128372 58108 128378 58172
rect 153326 58108 153332 58172
rect 153396 58108 153402 58172
rect 265198 58108 265204 58172
rect 265268 58108 265274 58172
rect 272190 58108 272196 58172
rect 272260 58108 272266 58172
rect 275686 58108 275692 58172
rect 275756 58108 275762 58172
rect 398230 58108 398236 58172
rect 398300 58108 398306 58172
rect 401726 58108 401732 58172
rect 401796 58108 401802 58172
rect 405406 58108 405412 58172
rect 405476 58108 405482 58172
rect 455822 58108 455828 58172
rect 455892 58108 455898 58172
rect 83958 57972 83964 58036
rect 84028 58034 84034 58036
rect 84193 58034 84259 58037
rect 84028 58032 84259 58034
rect 84028 57976 84198 58032
rect 84254 57976 84259 58032
rect 84028 57974 84259 57976
rect 84028 57972 84034 57974
rect 84193 57971 84259 57974
rect 85438 57901 85498 58108
rect 92246 57901 92306 58108
rect 99422 57901 99482 58108
rect 128310 57901 128370 58108
rect 153334 57901 153394 58108
rect 76005 57900 76071 57901
rect 78213 57900 78279 57901
rect 79501 57900 79567 57901
rect 76005 57896 76052 57900
rect 76116 57898 76122 57900
rect 76005 57840 76010 57896
rect 76005 57836 76052 57840
rect 76116 57838 76162 57898
rect 78213 57896 78260 57900
rect 78324 57898 78330 57900
rect 78213 57840 78218 57896
rect 76116 57836 76122 57838
rect 78213 57836 78260 57840
rect 78324 57838 78370 57898
rect 79501 57896 79548 57900
rect 79612 57898 79618 57900
rect 80053 57898 80119 57901
rect 81893 57900 81959 57901
rect 80462 57898 80468 57900
rect 79501 57840 79506 57896
rect 78324 57836 78330 57838
rect 79501 57836 79548 57840
rect 79612 57838 79658 57898
rect 80053 57896 80468 57898
rect 80053 57840 80058 57896
rect 80114 57840 80468 57896
rect 80053 57838 80468 57840
rect 79612 57836 79618 57838
rect 76005 57835 76071 57836
rect 78213 57835 78279 57836
rect 79501 57835 79567 57836
rect 80053 57835 80119 57838
rect 80462 57836 80468 57838
rect 80532 57836 80538 57900
rect 81893 57896 81940 57900
rect 82004 57898 82010 57900
rect 81893 57840 81898 57896
rect 81893 57836 81940 57840
rect 82004 57838 82050 57898
rect 85389 57896 85498 57901
rect 85389 57840 85394 57896
rect 85450 57840 85498 57896
rect 85389 57838 85498 57840
rect 86493 57900 86559 57901
rect 86493 57896 86540 57900
rect 86604 57898 86610 57900
rect 86953 57898 87019 57901
rect 88701 57900 88767 57901
rect 87638 57898 87644 57900
rect 86493 57840 86498 57896
rect 82004 57836 82010 57838
rect 81893 57835 81959 57836
rect 85389 57835 85455 57838
rect 86493 57836 86540 57840
rect 86604 57838 86650 57898
rect 86953 57896 87644 57898
rect 86953 57840 86958 57896
rect 87014 57840 87644 57896
rect 86953 57838 87644 57840
rect 86604 57836 86610 57838
rect 86493 57835 86559 57836
rect 86953 57835 87019 57838
rect 87638 57836 87644 57838
rect 87708 57836 87714 57900
rect 88701 57896 88748 57900
rect 88812 57898 88818 57900
rect 89805 57898 89871 57901
rect 90725 57900 90791 57901
rect 90030 57898 90036 57900
rect 88701 57840 88706 57896
rect 88701 57836 88748 57840
rect 88812 57838 88858 57898
rect 89805 57896 90036 57898
rect 89805 57840 89810 57896
rect 89866 57840 90036 57896
rect 89805 57838 90036 57840
rect 88812 57836 88818 57838
rect 88701 57835 88767 57836
rect 89805 57835 89871 57838
rect 90030 57836 90036 57838
rect 90100 57836 90106 57900
rect 90725 57896 90772 57900
rect 90836 57898 90842 57900
rect 91185 57898 91251 57901
rect 91318 57898 91324 57900
rect 90725 57840 90730 57896
rect 90725 57836 90772 57840
rect 90836 57838 90882 57898
rect 91185 57896 91324 57898
rect 91185 57840 91190 57896
rect 91246 57840 91324 57896
rect 91185 57838 91324 57840
rect 90836 57836 90842 57838
rect 90725 57835 90791 57836
rect 91185 57835 91251 57838
rect 91318 57836 91324 57838
rect 91388 57836 91394 57900
rect 92197 57896 92306 57901
rect 92197 57840 92202 57896
rect 92258 57840 92306 57896
rect 92197 57838 92306 57840
rect 92473 57898 92539 57901
rect 93342 57898 93348 57900
rect 92473 57896 93348 57898
rect 92473 57840 92478 57896
rect 92534 57840 93348 57896
rect 92473 57838 93348 57840
rect 92197 57835 92263 57838
rect 92473 57835 92539 57838
rect 93342 57836 93348 57838
rect 93412 57836 93418 57900
rect 93577 57898 93643 57901
rect 93710 57898 93716 57900
rect 93577 57896 93716 57898
rect 93577 57840 93582 57896
rect 93638 57840 93716 57896
rect 93577 57838 93716 57840
rect 93577 57835 93643 57838
rect 93710 57836 93716 57838
rect 93780 57836 93786 57900
rect 99373 57896 99482 57901
rect 99373 57840 99378 57896
rect 99434 57840 99482 57896
rect 99373 57838 99482 57840
rect 109493 57900 109559 57901
rect 112069 57900 112135 57901
rect 109493 57896 109540 57900
rect 109604 57898 109610 57900
rect 109493 57840 109498 57896
rect 99373 57835 99439 57838
rect 109493 57836 109540 57840
rect 109604 57838 109650 57898
rect 112069 57896 112116 57900
rect 112180 57898 112186 57900
rect 113817 57898 113883 57901
rect 115933 57900 115999 57901
rect 114318 57898 114324 57900
rect 112069 57840 112074 57896
rect 109604 57836 109610 57838
rect 112069 57836 112116 57840
rect 112180 57838 112226 57898
rect 113817 57896 114324 57898
rect 113817 57840 113822 57896
rect 113878 57840 114324 57896
rect 113817 57838 114324 57840
rect 112180 57836 112186 57838
rect 109493 57835 109559 57836
rect 112069 57835 112135 57836
rect 113817 57835 113883 57838
rect 114318 57836 114324 57838
rect 114388 57836 114394 57900
rect 115933 57896 115980 57900
rect 116044 57898 116050 57900
rect 116669 57898 116735 57901
rect 123477 57900 123543 57901
rect 125869 57900 125935 57901
rect 116894 57898 116900 57900
rect 115933 57840 115938 57896
rect 115933 57836 115980 57840
rect 116044 57838 116090 57898
rect 116669 57896 116900 57898
rect 116669 57840 116674 57896
rect 116730 57840 116900 57896
rect 116669 57838 116900 57840
rect 116044 57836 116050 57838
rect 115933 57835 115999 57836
rect 116669 57835 116735 57838
rect 116894 57836 116900 57838
rect 116964 57836 116970 57900
rect 123477 57896 123524 57900
rect 123588 57898 123594 57900
rect 123477 57840 123482 57896
rect 123477 57836 123524 57840
rect 123588 57838 123634 57898
rect 125869 57896 125916 57900
rect 125980 57898 125986 57900
rect 125869 57840 125874 57896
rect 123588 57836 123594 57838
rect 125869 57836 125916 57840
rect 125980 57838 126026 57898
rect 128310 57896 128419 57901
rect 128310 57840 128358 57896
rect 128414 57840 128419 57896
rect 128310 57838 128419 57840
rect 125980 57836 125986 57838
rect 123477 57835 123543 57836
rect 125869 57835 125935 57836
rect 128353 57835 128419 57838
rect 130837 57900 130903 57901
rect 133413 57900 133479 57901
rect 145557 57900 145623 57901
rect 130837 57896 130884 57900
rect 130948 57898 130954 57900
rect 130837 57840 130842 57896
rect 130837 57836 130884 57840
rect 130948 57838 130994 57898
rect 133413 57896 133460 57900
rect 133524 57898 133530 57900
rect 133413 57840 133418 57896
rect 130948 57836 130954 57838
rect 133413 57836 133460 57840
rect 133524 57838 133570 57898
rect 145557 57896 145604 57900
rect 145668 57898 145674 57900
rect 145557 57840 145562 57896
rect 133524 57836 133530 57838
rect 145557 57836 145604 57840
rect 145668 57838 145714 57898
rect 153285 57896 153394 57901
rect 153285 57840 153290 57896
rect 153346 57840 153394 57896
rect 153285 57838 153394 57840
rect 145668 57836 145674 57838
rect 130837 57835 130903 57836
rect 133413 57835 133479 57836
rect 145557 57835 145623 57836
rect 153285 57835 153351 57838
rect 183134 57836 183140 57900
rect 183204 57898 183210 57900
rect 183277 57898 183343 57901
rect 183204 57896 183343 57898
rect 183204 57840 183282 57896
rect 183338 57840 183343 57896
rect 183204 57838 183343 57840
rect 183204 57836 183210 57838
rect 183277 57835 183343 57838
rect 237373 57898 237439 57901
rect 239213 57900 239279 57901
rect 238150 57898 238156 57900
rect 237373 57896 238156 57898
rect 237373 57840 237378 57896
rect 237434 57840 238156 57896
rect 237373 57838 238156 57840
rect 237373 57835 237439 57838
rect 238150 57836 238156 57838
rect 238220 57836 238226 57900
rect 239213 57896 239260 57900
rect 239324 57898 239330 57900
rect 240133 57898 240199 57901
rect 241605 57900 241671 57901
rect 242893 57900 242959 57901
rect 240542 57898 240548 57900
rect 239213 57840 239218 57896
rect 239213 57836 239260 57840
rect 239324 57838 239370 57898
rect 240133 57896 240548 57898
rect 240133 57840 240138 57896
rect 240194 57840 240548 57896
rect 240133 57838 240548 57840
rect 239324 57836 239330 57838
rect 239213 57835 239279 57836
rect 240133 57835 240199 57838
rect 240542 57836 240548 57838
rect 240612 57836 240618 57900
rect 241605 57896 241652 57900
rect 241716 57898 241722 57900
rect 241605 57840 241610 57896
rect 241605 57836 241652 57840
rect 241716 57838 241762 57898
rect 242893 57896 242940 57900
rect 243004 57898 243010 57900
rect 242893 57840 242898 57896
rect 241716 57836 241722 57838
rect 242893 57836 242940 57840
rect 243004 57838 243050 57898
rect 243004 57836 243010 57838
rect 244222 57836 244228 57900
rect 244292 57898 244298 57900
rect 244365 57898 244431 57901
rect 244292 57896 244431 57898
rect 244292 57840 244370 57896
rect 244426 57840 244431 57896
rect 244292 57838 244431 57840
rect 244292 57836 244298 57838
rect 241605 57835 241671 57836
rect 242893 57835 242959 57836
rect 244365 57835 244431 57838
rect 245285 57900 245351 57901
rect 245285 57896 245332 57900
rect 245396 57898 245402 57900
rect 245653 57898 245719 57901
rect 247677 57900 247743 57901
rect 246430 57898 246436 57900
rect 245285 57840 245290 57896
rect 245285 57836 245332 57840
rect 245396 57838 245442 57898
rect 245653 57896 246436 57898
rect 245653 57840 245658 57896
rect 245714 57840 246436 57896
rect 245653 57838 246436 57840
rect 245396 57836 245402 57838
rect 245285 57835 245351 57836
rect 245653 57835 245719 57838
rect 246430 57836 246436 57838
rect 246500 57836 246506 57900
rect 247677 57896 247724 57900
rect 247788 57898 247794 57900
rect 248413 57898 248479 57901
rect 250069 57900 250135 57901
rect 248638 57898 248644 57900
rect 247677 57840 247682 57896
rect 247677 57836 247724 57840
rect 247788 57838 247834 57898
rect 248413 57896 248644 57898
rect 248413 57840 248418 57896
rect 248474 57840 248644 57896
rect 248413 57838 248644 57840
rect 247788 57836 247794 57838
rect 247677 57835 247743 57836
rect 248413 57835 248479 57838
rect 248638 57836 248644 57838
rect 248708 57836 248714 57900
rect 250069 57896 250116 57900
rect 250180 57898 250186 57900
rect 250989 57898 251055 57901
rect 255998 57898 256004 57900
rect 250069 57840 250074 57896
rect 250069 57836 250116 57840
rect 250180 57838 250226 57898
rect 250989 57896 256004 57898
rect 250989 57840 250994 57896
rect 251050 57840 256004 57896
rect 250989 57838 256004 57840
rect 250180 57836 250186 57838
rect 250069 57835 250135 57836
rect 250989 57835 251055 57838
rect 255998 57836 256004 57838
rect 256068 57836 256074 57900
rect 264973 57898 265039 57901
rect 265206 57898 265266 58108
rect 271045 57900 271111 57901
rect 270902 57898 270908 57900
rect 258030 57838 264162 57898
rect 183461 57764 183527 57765
rect 57830 57700 57836 57764
rect 57900 57762 57906 57764
rect 117998 57762 118004 57764
rect 57900 57702 118004 57762
rect 57900 57700 57906 57702
rect 117998 57700 118004 57702
rect 118068 57700 118074 57764
rect 183461 57760 183508 57764
rect 183572 57762 183578 57764
rect 183461 57704 183466 57760
rect 183461 57700 183508 57704
rect 183572 57702 183618 57762
rect 183572 57700 183578 57702
rect 205030 57700 205036 57764
rect 205100 57762 205106 57764
rect 258030 57762 258090 57838
rect 205100 57702 258090 57762
rect 258349 57764 258415 57765
rect 258349 57760 258396 57764
rect 258460 57762 258466 57764
rect 263593 57762 263659 57765
rect 263910 57762 263916 57764
rect 258349 57704 258354 57760
rect 205100 57700 205106 57702
rect 258349 57700 258396 57704
rect 258460 57702 258506 57762
rect 263593 57760 263916 57762
rect 263593 57704 263598 57760
rect 263654 57704 263916 57760
rect 263593 57702 263916 57704
rect 258460 57700 258466 57702
rect 183461 57699 183527 57700
rect 258349 57699 258415 57700
rect 263593 57699 263659 57702
rect 263910 57700 263916 57702
rect 263980 57700 263986 57764
rect 264102 57762 264162 57838
rect 264973 57896 265266 57898
rect 264973 57840 264978 57896
rect 265034 57840 265266 57896
rect 264973 57838 265266 57840
rect 265390 57838 270908 57898
rect 264973 57835 265039 57838
rect 265390 57762 265450 57838
rect 270902 57836 270908 57838
rect 270972 57836 270978 57900
rect 271045 57896 271092 57900
rect 271156 57898 271162 57900
rect 271873 57898 271939 57901
rect 272198 57898 272258 58108
rect 271045 57840 271050 57896
rect 271045 57836 271092 57840
rect 271156 57838 271202 57898
rect 271873 57896 272258 57898
rect 271873 57840 271878 57896
rect 271934 57840 272258 57896
rect 271873 57838 272258 57840
rect 273253 57900 273319 57901
rect 273253 57896 273300 57900
rect 273364 57898 273370 57900
rect 274633 57898 274699 57901
rect 275694 57898 275754 58108
rect 273253 57840 273258 57896
rect 271156 57836 271162 57838
rect 271045 57835 271111 57836
rect 271873 57835 271939 57838
rect 273253 57836 273300 57840
rect 273364 57838 273410 57898
rect 274633 57896 275754 57898
rect 274633 57840 274638 57896
rect 274694 57840 275754 57896
rect 274633 57838 275754 57840
rect 276933 57900 276999 57901
rect 276933 57896 276980 57900
rect 277044 57898 277050 57900
rect 287605 57898 287671 57901
rect 293309 57900 293375 57901
rect 295885 57900 295951 57901
rect 288198 57898 288204 57900
rect 276933 57840 276938 57896
rect 273364 57836 273370 57838
rect 273253 57835 273319 57836
rect 274633 57835 274699 57838
rect 276933 57836 276980 57840
rect 277044 57838 277090 57898
rect 287605 57896 288204 57898
rect 287605 57840 287610 57896
rect 287666 57840 288204 57896
rect 287605 57838 288204 57840
rect 277044 57836 277050 57838
rect 276933 57835 276999 57836
rect 287605 57835 287671 57838
rect 288198 57836 288204 57838
rect 288268 57836 288274 57900
rect 293309 57896 293356 57900
rect 293420 57898 293426 57900
rect 293309 57840 293314 57896
rect 293309 57836 293356 57840
rect 293420 57838 293466 57898
rect 295885 57896 295932 57900
rect 295996 57898 296002 57900
rect 298093 57898 298159 57901
rect 303429 57900 303495 57901
rect 305821 57900 305887 57901
rect 310973 57900 311039 57901
rect 313365 57900 313431 57901
rect 298502 57898 298508 57900
rect 295885 57840 295890 57896
rect 293420 57836 293426 57838
rect 295885 57836 295932 57840
rect 295996 57838 296042 57898
rect 298093 57896 298508 57898
rect 298093 57840 298098 57896
rect 298154 57840 298508 57896
rect 298093 57838 298508 57840
rect 295996 57836 296002 57838
rect 293309 57835 293375 57836
rect 295885 57835 295951 57836
rect 298093 57835 298159 57838
rect 298502 57836 298508 57838
rect 298572 57836 298578 57900
rect 303429 57896 303476 57900
rect 303540 57898 303546 57900
rect 303429 57840 303434 57896
rect 303429 57836 303476 57840
rect 303540 57838 303586 57898
rect 305821 57896 305868 57900
rect 305932 57898 305938 57900
rect 305821 57840 305826 57896
rect 303540 57836 303546 57838
rect 305821 57836 305868 57840
rect 305932 57838 305978 57898
rect 310973 57896 311020 57900
rect 311084 57898 311090 57900
rect 310973 57840 310978 57896
rect 305932 57836 305938 57838
rect 310973 57836 311020 57840
rect 311084 57838 311130 57898
rect 313365 57896 313412 57900
rect 313476 57898 313482 57900
rect 318241 57898 318307 57901
rect 323301 57900 323367 57901
rect 343173 57900 343239 57901
rect 343449 57900 343515 57901
rect 318374 57898 318380 57900
rect 313365 57840 313370 57896
rect 311084 57836 311090 57838
rect 313365 57836 313412 57840
rect 313476 57838 313522 57898
rect 318241 57896 318380 57898
rect 318241 57840 318246 57896
rect 318302 57840 318380 57896
rect 318241 57838 318380 57840
rect 313476 57836 313482 57838
rect 303429 57835 303495 57836
rect 305821 57835 305887 57836
rect 310973 57835 311039 57836
rect 313365 57835 313431 57836
rect 318241 57835 318307 57838
rect 318374 57836 318380 57838
rect 318444 57836 318450 57900
rect 323301 57896 323348 57900
rect 323412 57898 323418 57900
rect 343173 57898 343220 57900
rect 323301 57840 323306 57896
rect 323301 57836 323348 57840
rect 323412 57838 323458 57898
rect 343128 57896 343220 57898
rect 343128 57840 343178 57896
rect 343128 57838 343220 57840
rect 323412 57836 323418 57838
rect 343173 57836 343220 57838
rect 343284 57836 343290 57900
rect 343398 57898 343404 57900
rect 343358 57838 343404 57898
rect 343468 57896 343515 57900
rect 343510 57840 343515 57896
rect 343398 57836 343404 57838
rect 343468 57836 343515 57840
rect 323301 57835 323367 57836
rect 343173 57835 343239 57836
rect 343449 57835 343515 57836
rect 397453 57898 397519 57901
rect 398238 57898 398298 58108
rect 401734 57901 401794 58108
rect 397453 57896 398298 57898
rect 397453 57840 397458 57896
rect 397514 57840 398298 57896
rect 397453 57838 398298 57840
rect 399477 57900 399543 57901
rect 399477 57896 399524 57900
rect 399588 57898 399594 57900
rect 400213 57898 400279 57901
rect 400438 57898 400444 57900
rect 399477 57840 399482 57896
rect 397453 57835 397519 57838
rect 399477 57836 399524 57840
rect 399588 57838 399634 57898
rect 400213 57896 400444 57898
rect 400213 57840 400218 57896
rect 400274 57840 400444 57896
rect 400213 57838 400444 57840
rect 399588 57836 399594 57838
rect 399477 57835 399543 57836
rect 400213 57835 400279 57838
rect 400438 57836 400444 57838
rect 400508 57836 400514 57900
rect 401685 57896 401794 57901
rect 401685 57840 401690 57896
rect 401746 57840 401794 57896
rect 401685 57838 401794 57840
rect 404353 57898 404419 57901
rect 405414 57898 405474 58108
rect 404353 57896 405474 57898
rect 404353 57840 404358 57896
rect 404414 57840 405474 57896
rect 404353 57838 405474 57840
rect 405825 57898 405891 57901
rect 406510 57898 406516 57900
rect 405825 57896 406516 57898
rect 405825 57840 405830 57896
rect 405886 57840 406516 57896
rect 405825 57838 406516 57840
rect 401685 57835 401751 57838
rect 404353 57835 404419 57838
rect 405825 57835 405891 57838
rect 406510 57836 406516 57838
rect 406580 57836 406586 57900
rect 407205 57898 407271 57901
rect 408309 57900 408375 57901
rect 408677 57900 408743 57901
rect 407614 57898 407620 57900
rect 407205 57896 407620 57898
rect 407205 57840 407210 57896
rect 407266 57840 407620 57896
rect 407205 57838 407620 57840
rect 407205 57835 407271 57838
rect 407614 57836 407620 57838
rect 407684 57836 407690 57900
rect 408309 57896 408356 57900
rect 408420 57898 408426 57900
rect 408309 57840 408314 57896
rect 408309 57836 408356 57840
rect 408420 57838 408466 57898
rect 408677 57896 408724 57900
rect 408788 57898 408794 57900
rect 409873 57898 409939 57901
rect 410006 57898 410012 57900
rect 408677 57840 408682 57896
rect 408420 57836 408426 57838
rect 408677 57836 408724 57840
rect 408788 57838 408834 57898
rect 409873 57896 410012 57898
rect 409873 57840 409878 57896
rect 409934 57840 410012 57896
rect 409873 57838 410012 57840
rect 408788 57836 408794 57838
rect 408309 57835 408375 57836
rect 408677 57835 408743 57836
rect 409873 57835 409939 57838
rect 410006 57836 410012 57838
rect 410076 57836 410082 57900
rect 411345 57898 411411 57901
rect 415485 57900 415551 57901
rect 425237 57900 425303 57901
rect 426433 57900 426499 57901
rect 412398 57898 412404 57900
rect 411345 57896 412404 57898
rect 411345 57840 411350 57896
rect 411406 57840 412404 57896
rect 411345 57838 412404 57840
rect 411345 57835 411411 57838
rect 412398 57836 412404 57838
rect 412468 57836 412474 57900
rect 415485 57896 415532 57900
rect 415596 57898 415602 57900
rect 415485 57840 415490 57896
rect 415485 57836 415532 57840
rect 415596 57838 415642 57898
rect 425237 57896 425284 57900
rect 425348 57898 425354 57900
rect 426382 57898 426388 57900
rect 425237 57840 425242 57896
rect 415596 57836 415602 57838
rect 425237 57836 425284 57840
rect 425348 57838 425394 57898
rect 426342 57838 426388 57898
rect 426452 57896 426499 57900
rect 426494 57840 426499 57896
rect 425348 57836 425354 57838
rect 426382 57836 426388 57838
rect 426452 57836 426499 57840
rect 415485 57835 415551 57836
rect 425237 57835 425303 57836
rect 426433 57835 426499 57836
rect 428549 57900 428615 57901
rect 428549 57896 428596 57900
rect 428660 57898 428666 57900
rect 429193 57898 429259 57901
rect 429694 57898 429700 57900
rect 428549 57840 428554 57896
rect 428549 57836 428596 57840
rect 428660 57838 428706 57898
rect 429193 57896 429700 57898
rect 429193 57840 429198 57896
rect 429254 57840 429700 57896
rect 429193 57838 429700 57840
rect 428660 57836 428666 57838
rect 428549 57835 428615 57836
rect 429193 57835 429259 57838
rect 429694 57836 429700 57838
rect 429764 57836 429770 57900
rect 430573 57898 430639 57901
rect 432229 57900 432295 57901
rect 433517 57900 433583 57901
rect 434621 57900 434687 57901
rect 435909 57900 435975 57901
rect 431166 57898 431172 57900
rect 430573 57896 431172 57898
rect 430573 57840 430578 57896
rect 430634 57840 431172 57896
rect 430573 57838 431172 57840
rect 430573 57835 430639 57838
rect 431166 57836 431172 57838
rect 431236 57836 431242 57900
rect 432229 57896 432276 57900
rect 432340 57898 432346 57900
rect 432229 57840 432234 57896
rect 432229 57836 432276 57840
rect 432340 57838 432386 57898
rect 433517 57896 433564 57900
rect 433628 57898 433634 57900
rect 433517 57840 433522 57896
rect 432340 57836 432346 57838
rect 433517 57836 433564 57840
rect 433628 57838 433674 57898
rect 434621 57896 434668 57900
rect 434732 57898 434738 57900
rect 434621 57840 434626 57896
rect 433628 57836 433634 57838
rect 434621 57836 434668 57840
rect 434732 57838 434778 57898
rect 435909 57896 435956 57900
rect 436020 57898 436026 57900
rect 436369 57898 436435 57901
rect 438485 57900 438551 57901
rect 445845 57900 445911 57901
rect 436870 57898 436876 57900
rect 435909 57840 435914 57896
rect 434732 57836 434738 57838
rect 435909 57836 435956 57840
rect 436020 57838 436066 57898
rect 436369 57896 436876 57898
rect 436369 57840 436374 57896
rect 436430 57840 436876 57896
rect 436369 57838 436876 57840
rect 436020 57836 436026 57838
rect 432229 57835 432295 57836
rect 433517 57835 433583 57836
rect 434621 57835 434687 57836
rect 435909 57835 435975 57836
rect 436369 57835 436435 57838
rect 436870 57836 436876 57838
rect 436940 57836 436946 57900
rect 438485 57896 438532 57900
rect 438596 57898 438602 57900
rect 438485 57840 438490 57896
rect 438485 57836 438532 57840
rect 438596 57838 438642 57898
rect 445845 57896 445892 57900
rect 445956 57898 445962 57900
rect 455830 57898 455890 58108
rect 445845 57840 445850 57896
rect 438596 57836 438602 57838
rect 445845 57836 445892 57840
rect 445956 57838 446002 57898
rect 451230 57838 455890 57898
rect 460933 57900 460999 57901
rect 465901 57900 465967 57901
rect 470869 57900 470935 57901
rect 478413 57900 478479 57901
rect 485957 57900 486023 57901
rect 460933 57896 460980 57900
rect 461044 57898 461050 57900
rect 460933 57840 460938 57896
rect 445956 57836 445962 57838
rect 438485 57835 438551 57836
rect 445845 57835 445911 57836
rect 264102 57702 265450 57762
rect 266445 57762 266511 57765
rect 267590 57762 267596 57764
rect 266445 57760 267596 57762
rect 266445 57704 266450 57760
rect 266506 57704 267596 57760
rect 266445 57702 267596 57704
rect 266445 57699 266511 57702
rect 267590 57700 267596 57702
rect 267660 57700 267666 57764
rect 268469 57762 268535 57765
rect 268694 57762 268700 57764
rect 268469 57760 268700 57762
rect 268469 57704 268474 57760
rect 268530 57704 268700 57760
rect 268469 57702 268700 57704
rect 268469 57699 268535 57702
rect 268694 57700 268700 57702
rect 268764 57700 268770 57764
rect 269113 57762 269179 57765
rect 269798 57762 269804 57764
rect 269113 57760 269804 57762
rect 269113 57704 269118 57760
rect 269174 57704 269804 57760
rect 269113 57702 269804 57704
rect 269113 57699 269179 57702
rect 269798 57700 269804 57702
rect 269868 57700 269874 57764
rect 273345 57762 273411 57765
rect 274398 57762 274404 57764
rect 273345 57760 274404 57762
rect 273345 57704 273350 57760
rect 273406 57704 274404 57760
rect 273345 57702 274404 57704
rect 273345 57699 273411 57702
rect 274398 57700 274404 57702
rect 274468 57700 274474 57764
rect 358118 57700 358124 57764
rect 358188 57762 358194 57764
rect 443494 57762 443500 57764
rect 358188 57702 443500 57762
rect 358188 57700 358194 57702
rect 443494 57700 443500 57702
rect 443564 57700 443570 57764
rect 57646 57564 57652 57628
rect 57716 57626 57722 57628
rect 106273 57626 106339 57629
rect 106406 57626 106412 57628
rect 57716 57566 98746 57626
rect 57716 57564 57722 57566
rect 58566 57428 58572 57492
rect 58636 57490 58642 57492
rect 98545 57490 98611 57493
rect 58636 57488 98611 57490
rect 58636 57432 98550 57488
rect 98606 57432 98611 57488
rect 58636 57430 98611 57432
rect 98686 57490 98746 57566
rect 106273 57624 106412 57626
rect 106273 57568 106278 57624
rect 106334 57568 106412 57624
rect 106273 57566 106412 57568
rect 106273 57563 106339 57566
rect 106406 57564 106412 57566
rect 106476 57564 106482 57628
rect 110413 57626 110479 57629
rect 113265 57628 113331 57629
rect 111190 57626 111196 57628
rect 110413 57624 111196 57626
rect 110413 57568 110418 57624
rect 110474 57568 111196 57624
rect 110413 57566 111196 57568
rect 110413 57563 110479 57566
rect 111190 57564 111196 57566
rect 111260 57564 111266 57628
rect 113214 57626 113220 57628
rect 113174 57566 113220 57626
rect 113284 57624 113331 57628
rect 113326 57568 113331 57624
rect 113214 57564 113220 57566
rect 113284 57564 113331 57568
rect 113265 57563 113331 57564
rect 114553 57626 114619 57629
rect 115790 57626 115796 57628
rect 114553 57624 115796 57626
rect 114553 57568 114558 57624
rect 114614 57568 115796 57624
rect 114553 57566 115796 57568
rect 114553 57563 114619 57566
rect 115790 57564 115796 57566
rect 115860 57564 115866 57628
rect 118693 57626 118759 57629
rect 155953 57628 156019 57629
rect 119102 57626 119108 57628
rect 118693 57624 119108 57626
rect 118693 57568 118698 57624
rect 118754 57568 119108 57624
rect 118693 57566 119108 57568
rect 118693 57563 118759 57566
rect 119102 57564 119108 57566
rect 119172 57564 119178 57628
rect 155902 57626 155908 57628
rect 155862 57566 155908 57626
rect 155972 57624 156019 57628
rect 156014 57568 156019 57624
rect 155902 57564 155908 57566
rect 155972 57564 156019 57568
rect 155953 57563 156019 57564
rect 160093 57626 160159 57629
rect 160870 57626 160876 57628
rect 160093 57624 160876 57626
rect 160093 57568 160098 57624
rect 160154 57568 160876 57624
rect 160093 57566 160876 57568
rect 160093 57563 160159 57566
rect 160870 57564 160876 57566
rect 160940 57564 160946 57628
rect 165613 57626 165679 57629
rect 165838 57626 165844 57628
rect 165613 57624 165844 57626
rect 165613 57568 165618 57624
rect 165674 57568 165844 57624
rect 165613 57566 165844 57568
rect 165613 57563 165679 57566
rect 165838 57564 165844 57566
rect 165908 57564 165914 57628
rect 213126 57564 213132 57628
rect 213196 57626 213202 57628
rect 278446 57626 278452 57628
rect 213196 57566 278452 57626
rect 213196 57564 213202 57566
rect 278446 57564 278452 57566
rect 278516 57564 278522 57628
rect 374678 57564 374684 57628
rect 374748 57626 374754 57628
rect 451230 57626 451290 57838
rect 460933 57836 460980 57840
rect 461044 57838 461090 57898
rect 465901 57896 465948 57900
rect 466012 57898 466018 57900
rect 465901 57840 465906 57896
rect 461044 57836 461050 57838
rect 465901 57836 465948 57840
rect 466012 57838 466058 57898
rect 470869 57896 470916 57900
rect 470980 57898 470986 57900
rect 470869 57840 470874 57896
rect 466012 57836 466018 57838
rect 470869 57836 470916 57840
rect 470980 57838 471026 57898
rect 478413 57896 478460 57900
rect 478524 57898 478530 57900
rect 478413 57840 478418 57896
rect 470980 57836 470986 57838
rect 478413 57836 478460 57840
rect 478524 57838 478570 57898
rect 485957 57896 486004 57900
rect 486068 57898 486074 57900
rect 485957 57840 485962 57896
rect 478524 57836 478530 57838
rect 485957 57836 486004 57840
rect 486068 57838 486114 57898
rect 486068 57836 486074 57838
rect 503110 57836 503116 57900
rect 503180 57898 503186 57900
rect 503253 57898 503319 57901
rect 503529 57900 503595 57901
rect 503180 57896 503319 57898
rect 503180 57840 503258 57896
rect 503314 57840 503319 57896
rect 503180 57838 503319 57840
rect 503180 57836 503186 57838
rect 460933 57835 460999 57836
rect 465901 57835 465967 57836
rect 470869 57835 470935 57836
rect 478413 57835 478479 57836
rect 485957 57835 486023 57836
rect 503253 57835 503319 57838
rect 503478 57836 503484 57900
rect 503548 57898 503595 57900
rect 503548 57896 503640 57898
rect 503590 57840 503640 57896
rect 503548 57838 503640 57840
rect 503548 57836 503595 57838
rect 503529 57835 503595 57836
rect 374748 57566 451290 57626
rect 374748 57564 374754 57566
rect 105302 57490 105308 57492
rect 98686 57430 105308 57490
rect 58636 57428 58642 57430
rect 98545 57427 98611 57430
rect 105302 57428 105308 57430
rect 105372 57428 105378 57492
rect 203190 57428 203196 57492
rect 203260 57490 203266 57492
rect 250989 57490 251055 57493
rect 203260 57488 251055 57490
rect 203260 57432 250994 57488
rect 251050 57432 251055 57488
rect 203260 57430 251055 57432
rect 203260 57428 203266 57430
rect 250989 57427 251055 57430
rect 251173 57492 251239 57493
rect 251173 57488 251220 57492
rect 251284 57490 251290 57492
rect 251909 57490 251975 57493
rect 252318 57490 252324 57492
rect 251173 57432 251178 57488
rect 251173 57428 251220 57432
rect 251284 57430 251330 57490
rect 251909 57488 252324 57490
rect 251909 57432 251914 57488
rect 251970 57432 252324 57488
rect 251909 57430 252324 57432
rect 251284 57428 251290 57430
rect 251173 57427 251239 57428
rect 251909 57427 251975 57430
rect 252318 57428 252324 57430
rect 252388 57428 252394 57492
rect 252553 57490 252619 57493
rect 253422 57490 253428 57492
rect 252553 57488 253428 57490
rect 252553 57432 252558 57488
rect 252614 57432 253428 57488
rect 252553 57430 253428 57432
rect 252553 57427 252619 57430
rect 253422 57428 253428 57430
rect 253492 57428 253498 57492
rect 253933 57490 253999 57493
rect 266353 57492 266419 57493
rect 254526 57490 254532 57492
rect 253933 57488 254532 57490
rect 253933 57432 253938 57488
rect 253994 57432 254532 57488
rect 253933 57430 254532 57432
rect 253933 57427 253999 57430
rect 254526 57428 254532 57430
rect 254596 57428 254602 57492
rect 266302 57490 266308 57492
rect 266262 57430 266308 57490
rect 266372 57488 266419 57492
rect 266414 57432 266419 57488
rect 266302 57428 266308 57430
rect 266372 57428 266419 57432
rect 370446 57428 370452 57492
rect 370516 57490 370522 57492
rect 433149 57490 433215 57493
rect 433425 57492 433491 57493
rect 433374 57490 433380 57492
rect 370516 57488 433215 57490
rect 370516 57432 433154 57488
rect 433210 57432 433215 57488
rect 370516 57430 433215 57432
rect 433334 57430 433380 57490
rect 433444 57488 433491 57492
rect 433486 57432 433491 57488
rect 370516 57428 370522 57430
rect 266353 57427 266419 57428
rect 433149 57427 433215 57430
rect 433374 57428 433380 57430
rect 433444 57428 433491 57432
rect 433425 57427 433491 57428
rect 434713 57490 434779 57493
rect 435766 57490 435772 57492
rect 434713 57488 435772 57490
rect 434713 57432 434718 57488
rect 434774 57432 435772 57488
rect 434713 57430 435772 57432
rect 434713 57427 434779 57430
rect 435766 57428 435772 57430
rect 435836 57428 435842 57492
rect 437473 57490 437539 57493
rect 438342 57490 438348 57492
rect 437473 57488 438348 57490
rect 437473 57432 437478 57488
rect 437534 57432 438348 57488
rect 437473 57430 438348 57432
rect 437473 57427 437539 57430
rect 438342 57428 438348 57430
rect 438412 57428 438418 57492
rect 58750 57292 58756 57356
rect 58820 57354 58826 57356
rect 98494 57354 98500 57356
rect 58820 57294 98500 57354
rect 58820 57292 58826 57294
rect 98494 57292 98500 57294
rect 98564 57292 98570 57356
rect 213310 57292 213316 57356
rect 213380 57354 213386 57356
rect 265934 57354 265940 57356
rect 213380 57294 265940 57354
rect 213380 57292 213386 57294
rect 265934 57292 265940 57294
rect 266004 57292 266010 57356
rect 379094 57292 379100 57356
rect 379164 57354 379170 57356
rect 448278 57354 448284 57356
rect 379164 57294 448284 57354
rect 379164 57292 379170 57294
rect 448278 57292 448284 57294
rect 448348 57292 448354 57356
rect 50470 57156 50476 57220
rect 50540 57218 50546 57220
rect 88374 57218 88380 57220
rect 50540 57158 88380 57218
rect 50540 57156 50546 57158
rect 88374 57156 88380 57158
rect 88444 57156 88450 57220
rect 98545 57218 98611 57221
rect 103830 57218 103836 57220
rect 98545 57216 103836 57218
rect 98545 57160 98550 57216
rect 98606 57160 103836 57216
rect 98545 57158 103836 57160
rect 98545 57155 98611 57158
rect 103830 57156 103836 57158
rect 103900 57156 103906 57220
rect 202086 57156 202092 57220
rect 202156 57218 202162 57220
rect 248270 57218 248276 57220
rect 202156 57158 248276 57218
rect 202156 57156 202162 57158
rect 248270 57156 248276 57158
rect 248340 57156 248346 57220
rect 378910 57156 378916 57220
rect 378980 57218 378986 57220
rect 418470 57218 418476 57220
rect 378980 57158 418476 57218
rect 378980 57156 378986 57158
rect 418470 57156 418476 57158
rect 418540 57156 418546 57220
rect 426525 57218 426591 57221
rect 430941 57220 431007 57221
rect 427670 57218 427676 57220
rect 426525 57216 427676 57218
rect 426525 57160 426530 57216
rect 426586 57160 427676 57216
rect 426525 57158 427676 57160
rect 426525 57155 426591 57158
rect 427670 57156 427676 57158
rect 427740 57156 427746 57220
rect 430941 57216 430988 57220
rect 431052 57218 431058 57220
rect 433149 57218 433215 57221
rect 440918 57218 440924 57220
rect 430941 57160 430946 57216
rect 430941 57156 430988 57160
rect 431052 57158 431098 57218
rect 433149 57216 440924 57218
rect 433149 57160 433154 57216
rect 433210 57160 440924 57216
rect 433149 57158 440924 57160
rect 431052 57156 431058 57158
rect 430941 57155 431007 57156
rect 433149 57155 433215 57158
rect 440918 57156 440924 57158
rect 440988 57156 440994 57220
rect 58934 57020 58940 57084
rect 59004 57082 59010 57084
rect 96286 57082 96292 57084
rect 59004 57022 96292 57082
rect 59004 57020 59010 57022
rect 96286 57020 96292 57022
rect 96356 57020 96362 57084
rect 215886 57020 215892 57084
rect 215956 57082 215962 57084
rect 260966 57082 260972 57084
rect 215956 57022 260972 57082
rect 215956 57020 215962 57022
rect 260966 57020 260972 57022
rect 261036 57020 261042 57084
rect 378726 57020 378732 57084
rect 378796 57082 378802 57084
rect 413502 57082 413508 57084
rect 378796 57022 413508 57082
rect 378796 57020 378802 57022
rect 413502 57020 413508 57022
rect 413572 57020 413578 57084
rect 411253 56948 411319 56949
rect 411253 56944 411300 56948
rect 411364 56946 411370 56948
rect 412541 56946 412607 56949
rect 411253 56888 411258 56944
rect 411253 56884 411300 56888
rect 411364 56886 411410 56946
rect 412541 56944 412650 56946
rect 412541 56888 412546 56944
rect 412602 56888 412650 56944
rect 411364 56884 411370 56886
rect 411253 56883 411319 56884
rect 412541 56883 412650 56888
rect 412590 56813 412650 56883
rect 55070 56748 55076 56812
rect 55140 56810 55146 56812
rect 118366 56810 118372 56812
rect 55140 56750 118372 56810
rect 55140 56748 55146 56750
rect 118366 56748 118372 56750
rect 118436 56748 118442 56812
rect 412590 56808 412699 56813
rect 412590 56752 412638 56808
rect 412694 56752 412699 56808
rect 412590 56750 412699 56752
rect 412633 56747 412699 56750
rect 163262 56612 163268 56676
rect 163332 56612 163338 56676
rect 216070 56612 216076 56676
rect 216140 56674 216146 56676
rect 283782 56674 283788 56676
rect 216140 56614 283788 56674
rect 216140 56612 216146 56614
rect 283782 56612 283788 56614
rect 283852 56612 283858 56676
rect 360694 56612 360700 56676
rect 360764 56674 360770 56676
rect 451038 56674 451044 56676
rect 360764 56614 451044 56674
rect 360764 56612 360770 56614
rect 451038 56612 451044 56614
rect 451108 56612 451114 56676
rect 53598 56476 53604 56540
rect 53668 56538 53674 56540
rect 163270 56538 163330 56612
rect 53668 56478 163330 56538
rect 53668 56476 53674 56478
rect 219198 56476 219204 56540
rect 219268 56538 219274 56540
rect 426014 56538 426020 56540
rect 219268 56478 426020 56538
rect 219268 56476 219274 56478
rect 426014 56476 426020 56478
rect 426084 56476 426090 56540
rect 50654 56340 50660 56404
rect 50724 56402 50730 56404
rect 158478 56402 158484 56404
rect 50724 56342 158484 56402
rect 50724 56340 50730 56342
rect 158478 56340 158484 56342
rect 158548 56340 158554 56404
rect 219934 56340 219940 56404
rect 220004 56402 220010 56404
rect 421046 56402 421052 56404
rect 220004 56342 421052 56402
rect 220004 56340 220010 56342
rect 421046 56340 421052 56342
rect 421116 56340 421122 56404
rect 55622 56204 55628 56268
rect 55692 56266 55698 56268
rect 153285 56266 153351 56269
rect 55692 56264 153351 56266
rect 55692 56208 153290 56264
rect 153346 56208 153351 56264
rect 55692 56206 153351 56208
rect 55692 56204 55698 56206
rect 153285 56203 153351 56206
rect 201350 56204 201356 56268
rect 201420 56266 201426 56268
rect 273478 56266 273484 56268
rect 201420 56206 273484 56266
rect 201420 56204 201426 56206
rect 273478 56204 273484 56206
rect 273548 56204 273554 56268
rect 377622 56204 377628 56268
rect 377692 56266 377698 56268
rect 439078 56266 439084 56268
rect 377692 56206 439084 56266
rect 377692 56204 377698 56206
rect 439078 56204 439084 56206
rect 439148 56204 439154 56268
rect 217358 56068 217364 56132
rect 217428 56130 217434 56132
rect 277158 56130 277164 56132
rect 217428 56070 277164 56130
rect 217428 56068 217434 56070
rect 277158 56068 277164 56070
rect 277228 56068 277234 56132
rect 379462 56068 379468 56132
rect 379532 56130 379538 56132
rect 428549 56130 428615 56133
rect 379532 56128 428615 56130
rect 379532 56072 428554 56128
rect 428610 56072 428615 56128
rect 379532 56070 428615 56072
rect 379532 56068 379538 56070
rect 428549 56067 428615 56070
rect 377806 55932 377812 55996
rect 377876 55994 377882 55996
rect 425237 55994 425303 55997
rect 377876 55992 425303 55994
rect 377876 55936 425242 55992
rect 425298 55936 425303 55992
rect 377876 55934 425303 55936
rect 377876 55932 377882 55934
rect 425237 55931 425303 55934
rect 48630 55116 48636 55180
rect 48700 55178 48706 55180
rect 165613 55178 165679 55181
rect 48700 55176 165679 55178
rect 48700 55120 165618 55176
rect 165674 55120 165679 55176
rect 48700 55118 165679 55120
rect 48700 55116 48706 55118
rect 165613 55115 165679 55118
rect 213729 55178 213795 55181
rect 274633 55178 274699 55181
rect 213729 55176 274699 55178
rect 213729 55120 213734 55176
rect 213790 55120 274638 55176
rect 274694 55120 274699 55176
rect 213729 55118 274699 55120
rect 213729 55115 213795 55118
rect 274633 55115 274699 55118
rect 50838 54980 50844 55044
rect 50908 55042 50914 55044
rect 160093 55042 160159 55045
rect 50908 55040 160159 55042
rect 50908 54984 160098 55040
rect 160154 54984 160159 55040
rect 50908 54982 160159 54984
rect 50908 54980 50914 54982
rect 160093 54979 160159 54982
rect 214925 55042 214991 55045
rect 269113 55042 269179 55045
rect 214925 55040 269179 55042
rect 214925 54984 214930 55040
rect 214986 54984 269118 55040
rect 269174 54984 269179 55040
rect 214925 54982 269179 54984
rect 214925 54979 214991 54982
rect 269113 54979 269179 54982
rect 52310 54844 52316 54908
rect 52380 54906 52386 54908
rect 155953 54906 156019 54909
rect 52380 54904 156019 54906
rect 52380 54848 155958 54904
rect 156014 54848 156019 54904
rect 52380 54846 156019 54848
rect 52380 54844 52386 54846
rect 155953 54843 156019 54846
rect 57462 54708 57468 54772
rect 57532 54770 57538 54772
rect 118693 54770 118759 54773
rect 57532 54768 118759 54770
rect 57532 54712 118698 54768
rect 118754 54712 118759 54768
rect 57532 54710 118759 54712
rect 57532 54708 57538 54710
rect 118693 54707 118759 54710
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 136449 4042 136515 4045
rect 204846 4042 204852 4044
rect 136449 4040 204852 4042
rect 136449 3984 136454 4040
rect 136510 3984 204852 4040
rect 136449 3982 204852 3984
rect 136449 3979 136515 3982
rect 204846 3980 204852 3982
rect 204916 3980 204922 4044
rect 140037 3906 140103 3909
rect 210366 3906 210372 3908
rect 140037 3904 210372 3906
rect 140037 3848 140042 3904
rect 140098 3848 210372 3904
rect 140037 3846 210372 3848
rect 140037 3843 140103 3846
rect 210366 3844 210372 3846
rect 210436 3844 210442 3908
rect 147121 3770 147187 3773
rect 363454 3770 363460 3772
rect 147121 3768 363460 3770
rect 147121 3712 147126 3768
rect 147182 3712 363460 3768
rect 147121 3710 363460 3712
rect 147121 3707 147187 3710
rect 363454 3708 363460 3710
rect 363524 3708 363530 3772
rect 150617 3634 150683 3637
rect 367870 3634 367876 3636
rect 150617 3632 367876 3634
rect 150617 3576 150622 3632
rect 150678 3576 367876 3632
rect 150617 3574 367876 3576
rect 150617 3571 150683 3574
rect 367870 3572 367876 3574
rect 367940 3572 367946 3636
rect 132953 3498 133019 3501
rect 363638 3498 363644 3500
rect 132953 3496 363644 3498
rect 132953 3440 132958 3496
rect 133014 3440 363644 3496
rect 132953 3438 363644 3440
rect 132953 3435 133019 3438
rect 363638 3436 363644 3438
rect 363708 3436 363714 3500
rect 129365 3362 129431 3365
rect 367686 3362 367692 3364
rect 129365 3360 367692 3362
rect 129365 3304 129370 3360
rect 129426 3304 367692 3360
rect 129365 3302 367692 3304
rect 129365 3299 129431 3302
rect 367686 3300 367692 3302
rect 367756 3300 367762 3364
rect 143533 3226 143599 3229
rect 206134 3226 206140 3228
rect 143533 3224 206140 3226
rect 143533 3168 143538 3224
rect 143594 3168 206140 3224
rect 143533 3166 206140 3168
rect 143533 3163 143599 3166
rect 206134 3164 206140 3166
rect 206204 3164 206210 3228
<< via3 >>
rect 54340 632572 54404 632636
rect 53052 632436 53116 632500
rect 476068 627812 476132 627876
rect 488580 627812 488644 627876
rect 506612 627812 506676 627876
rect 121684 618428 121748 618492
rect 436140 594764 436204 594828
rect 121684 552604 121748 552668
rect 299980 549476 300044 549540
rect 299980 522548 300044 522612
rect 436140 522276 436204 522340
rect 360884 516700 360948 516764
rect 363460 515340 363524 515404
rect 363644 491812 363708 491876
rect 476068 491812 476132 491876
rect 367692 490452 367756 490516
rect 367876 487732 367940 487796
rect 206140 486372 206204 486436
rect 488580 486372 488644 486436
rect 59308 485692 59372 485756
rect 196756 485692 196820 485756
rect 212396 485692 212460 485756
rect 357940 485692 358004 485756
rect 54708 485556 54772 485620
rect 202276 485556 202340 485620
rect 213684 485556 213748 485620
rect 364932 485556 364996 485620
rect 51948 485420 52012 485484
rect 196572 485420 196636 485484
rect 371740 485420 371804 485484
rect 53420 485284 53484 485348
rect 197860 485284 197924 485348
rect 217548 485284 217612 485348
rect 373764 485284 373828 485348
rect 50292 485148 50356 485212
rect 198596 485148 198660 485212
rect 205404 485148 205468 485212
rect 206876 485148 206940 485212
rect 219204 485148 219268 485212
rect 374500 485148 374564 485212
rect 57836 485012 57900 485076
rect 200620 485012 200684 485076
rect 208900 485012 208964 485076
rect 219020 485012 219084 485076
rect 375972 485012 376036 485076
rect 59124 484876 59188 484940
rect 198044 484876 198108 484940
rect 202644 484876 202708 484940
rect 356652 484876 356716 484940
rect 198412 484740 198476 484804
rect 201356 484740 201420 484804
rect 209084 484740 209148 484804
rect 200804 484604 200868 484668
rect 211660 484604 211724 484668
rect 53236 484528 53300 484532
rect 53236 484472 53286 484528
rect 53286 484472 53300 484528
rect 53236 484468 53300 484472
rect 53604 484528 53668 484532
rect 53604 484472 53654 484528
rect 53654 484472 53668 484528
rect 53604 484468 53668 484472
rect 216996 484468 217060 484532
rect 219940 484468 220004 484532
rect 377444 483924 377508 483988
rect 205772 483788 205836 483852
rect 377260 483788 377324 483852
rect 213132 483652 213196 483716
rect 360700 483652 360764 483716
rect 46796 482836 46860 482900
rect 47716 482700 47780 482764
rect 375420 482428 375484 482492
rect 213868 482292 213932 482356
rect 376156 482292 376220 482356
rect 215340 480932 215404 480996
rect 374868 480932 374932 480996
rect 215892 480796 215956 480860
rect 370084 480796 370148 480860
rect 57468 479844 57532 479908
rect 57100 479708 57164 479772
rect 217180 479708 217244 479772
rect 44956 479572 45020 479636
rect 213316 479572 213380 479636
rect 364380 479572 364444 479636
rect 44772 479436 44836 479500
rect 208348 479436 208412 479500
rect 210372 479436 210436 479500
rect 209820 478212 209884 478276
rect 378732 478212 378796 478276
rect 198964 478076 199028 478140
rect 204852 478076 204916 478140
rect 376892 476988 376956 477052
rect 203196 476852 203260 476916
rect 370452 476852 370516 476916
rect 214052 476716 214116 476780
rect 378180 476716 378244 476780
rect 210004 475492 210068 475556
rect 377628 475492 377692 475556
rect 216076 475356 216140 475420
rect 359412 475356 359476 475420
rect 359780 474540 359844 474604
rect 358124 474404 358188 474468
rect 379468 474268 379532 474332
rect 374684 474132 374748 474196
rect 214420 473996 214484 474060
rect 378916 473996 378980 474060
rect 205220 472772 205284 472836
rect 206324 472636 206388 472700
rect 506612 472636 506676 472700
rect 202092 472500 202156 472564
rect 379100 472500 379164 472564
rect 202460 471684 202524 471748
rect 207980 471548 208044 471612
rect 47900 471412 47964 471476
rect 217364 471412 217428 471476
rect 214604 471140 214668 471204
rect 58940 469780 59004 469844
rect 205036 469780 205100 469844
rect 58756 469100 58820 469164
rect 199516 469100 199580 469164
rect 48084 468964 48148 469028
rect 200988 468964 201052 469028
rect 52316 468828 52380 468892
rect 203012 468828 203076 468892
rect 50844 468692 50908 468756
rect 50660 468556 50724 468620
rect 213500 468556 213564 468620
rect 48636 468420 48700 468484
rect 208164 468420 208228 468484
rect 359596 468420 359660 468484
rect 60228 467196 60292 467260
rect 179644 467196 179708 467260
rect 44036 467060 44100 467124
rect 218652 467060 218716 467124
rect 359964 467060 360028 467124
rect 178356 466516 178420 466580
rect 190868 466576 190932 466580
rect 190868 466520 190918 466576
rect 190918 466520 190932 466576
rect 190868 466516 190932 466520
rect 338436 466576 338500 466580
rect 338436 466520 338486 466576
rect 338486 466520 338500 466576
rect 338436 466516 338500 466520
rect 339724 466576 339788 466580
rect 339724 466520 339774 466576
rect 339774 466520 339788 466576
rect 339724 466516 339788 466520
rect 350948 466576 351012 466580
rect 350948 466520 350998 466576
rect 350998 466520 351012 466576
rect 350948 466516 351012 466520
rect 498516 466576 498580 466580
rect 498516 466520 498530 466576
rect 498530 466520 498580 466576
rect 498516 466516 498580 466520
rect 499804 466576 499868 466580
rect 499804 466520 499818 466576
rect 499818 466520 499868 466576
rect 499804 466516 499868 466520
rect 510844 466576 510908 466580
rect 510844 466520 510894 466576
rect 510894 466520 510908 466576
rect 510844 466516 510908 466520
rect 50476 466380 50540 466444
rect 55076 466244 55140 466308
rect 198780 466244 198844 466308
rect 55444 466108 55508 466172
rect 54892 465972 54956 466036
rect 46612 465836 46676 465900
rect 52132 465700 52196 465764
rect 58572 465564 58636 465628
rect 51580 465156 51644 465220
rect 55628 465216 55692 465220
rect 55628 465160 55678 465216
rect 55678 465160 55692 465216
rect 55628 465156 55692 465160
rect 199148 464340 199212 464404
rect 205404 411300 205468 411364
rect 199148 397972 199212 398036
rect 199148 396128 199212 396132
rect 199148 396072 199198 396128
rect 199198 396072 199212 396128
rect 199148 396068 199212 396072
rect 199332 395796 199396 395860
rect 208348 390628 208412 390692
rect 51948 388452 52012 388516
rect 57652 388452 57716 388516
rect 377628 382332 377692 382396
rect 359964 381516 360028 381580
rect 59860 380972 59924 381036
rect 205588 380972 205652 381036
rect 93462 380836 93526 380900
rect 111006 380896 111070 380900
rect 111006 380840 111026 380896
rect 111026 380840 111070 380896
rect 111006 380836 111070 380840
rect 113590 380896 113654 380900
rect 113590 380840 113602 380896
rect 113602 380840 113654 380896
rect 113590 380836 113654 380840
rect 116038 380896 116102 380900
rect 116038 380840 116086 380896
rect 116086 380840 116102 380896
rect 116038 380836 116102 380840
rect 118486 380836 118550 380900
rect 120934 380836 120998 380900
rect 123518 380896 123582 380900
rect 123518 380840 123538 380896
rect 123538 380840 123582 380896
rect 123518 380836 123582 380840
rect 125966 380896 126030 380900
rect 125966 380840 126022 380896
rect 126022 380840 126030 380896
rect 125966 380836 126030 380840
rect 130998 380896 131062 380900
rect 130998 380840 131026 380896
rect 131026 380840 131062 380896
rect 130998 380836 131062 380840
rect 133446 380836 133510 380900
rect 135894 380896 135958 380900
rect 135894 380840 135902 380896
rect 135902 380840 135958 380896
rect 135894 380836 135958 380840
rect 143510 380896 143574 380900
rect 143510 380840 143538 380896
rect 143538 380840 143574 380896
rect 143510 380836 143574 380840
rect 145958 380836 146022 380900
rect 158470 380836 158534 380900
rect 160918 380896 160982 380900
rect 160918 380840 160926 380896
rect 160926 380840 160982 380896
rect 160918 380836 160982 380840
rect 163366 380896 163430 380900
rect 163366 380840 163410 380896
rect 163410 380840 163430 380896
rect 163366 380836 163430 380840
rect 165950 380896 166014 380900
rect 165950 380840 165986 380896
rect 165986 380840 166014 380896
rect 165950 380836 166014 380840
rect 263934 380836 263998 380900
rect 485950 380836 486014 380900
rect 236054 380700 236118 380764
rect 237142 380760 237206 380764
rect 237142 380704 237158 380760
rect 237158 380704 237206 380760
rect 237142 380700 237206 380704
rect 243126 380760 243190 380764
rect 243126 380704 243138 380760
rect 243138 380704 243190 380760
rect 243126 380700 243190 380704
rect 245438 380700 245502 380764
rect 256046 380760 256110 380764
rect 256046 380704 256054 380760
rect 256054 380704 256110 380760
rect 256046 380700 256110 380704
rect 269782 380760 269846 380764
rect 269782 380704 269818 380760
rect 269818 380704 269846 380760
rect 269782 380700 269846 380704
rect 421078 380760 421142 380764
rect 421078 380704 421102 380760
rect 421102 380704 421142 380760
rect 421078 380700 421142 380704
rect 422846 380760 422910 380764
rect 422846 380704 422850 380760
rect 422850 380704 422906 380760
rect 422906 380704 422910 380760
rect 422846 380700 422910 380704
rect 431006 380700 431070 380764
rect 433590 380760 433654 380764
rect 433590 380704 433614 380760
rect 433614 380704 433654 380760
rect 433590 380700 433654 380704
rect 436038 380760 436102 380764
rect 436038 380704 436062 380760
rect 436062 380704 436102 380760
rect 436038 380700 436102 380704
rect 438486 380760 438550 380764
rect 438486 380704 438490 380760
rect 438490 380704 438546 380760
rect 438546 380704 438550 380760
rect 438486 380700 438550 380704
rect 440934 380760 440998 380764
rect 440934 380704 440938 380760
rect 440938 380704 440998 380760
rect 440934 380700 440998 380704
rect 443518 380700 443582 380764
rect 77142 380564 77206 380628
rect 76052 380428 76116 380492
rect 128308 380352 128372 380356
rect 128308 380296 128358 380352
rect 128358 380296 128372 380352
rect 128308 380292 128372 380296
rect 155908 380352 155972 380356
rect 155908 380296 155958 380352
rect 155958 380296 155972 380352
rect 155908 380292 155972 380296
rect 216628 380428 216692 380492
rect 216996 380428 217060 380492
rect 254550 380564 254614 380628
rect 255910 380624 255974 380628
rect 255910 380568 255926 380624
rect 255926 380568 255974 380624
rect 255910 380564 255974 380568
rect 256998 380624 257062 380628
rect 256998 380568 257030 380624
rect 257030 380568 257062 380624
rect 256998 380564 257062 380568
rect 259446 380624 259510 380628
rect 259446 380568 259458 380624
rect 259458 380568 259510 380624
rect 259446 380564 259510 380568
rect 260670 380564 260734 380628
rect 265294 380624 265358 380628
rect 265294 380568 265310 380624
rect 265310 380568 265358 380624
rect 265294 380564 265358 380568
rect 271006 380624 271070 380628
rect 271006 380568 271014 380624
rect 271014 380568 271070 380624
rect 271006 380564 271070 380568
rect 408702 380624 408766 380628
rect 408702 380568 408738 380624
rect 408738 380568 408766 380624
rect 408702 380564 408766 380568
rect 413462 380624 413526 380628
rect 413462 380568 413466 380624
rect 413466 380568 413522 380624
rect 413522 380568 413526 380624
rect 413462 380564 413526 380568
rect 419446 380624 419510 380628
rect 419446 380568 419502 380624
rect 419502 380568 419510 380624
rect 419446 380564 419510 380568
rect 434406 380564 434470 380628
rect 445966 380624 446030 380628
rect 445966 380568 445998 380624
rect 445998 380568 446030 380624
rect 445966 380564 446030 380568
rect 119108 380156 119172 380220
rect 50292 379476 50356 379540
rect 202644 379476 202708 379540
rect 209084 379476 209148 379540
rect 364380 379476 364444 379540
rect 79548 379340 79612 379404
rect 85436 379400 85500 379404
rect 85436 379344 85486 379400
rect 85486 379344 85500 379400
rect 85436 379340 85500 379344
rect 86540 379400 86604 379404
rect 86540 379344 86590 379400
rect 86590 379344 86604 379400
rect 86540 379340 86604 379344
rect 87644 379400 87708 379404
rect 87644 379344 87694 379400
rect 87694 379344 87708 379400
rect 87644 379340 87708 379344
rect 88380 379400 88444 379404
rect 88380 379344 88394 379400
rect 88394 379344 88444 379400
rect 88380 379340 88444 379344
rect 88748 379400 88812 379404
rect 88748 379344 88798 379400
rect 88798 379344 88812 379400
rect 88748 379340 88812 379344
rect 90036 379400 90100 379404
rect 90036 379344 90086 379400
rect 90086 379344 90100 379400
rect 90036 379340 90100 379344
rect 90772 379340 90836 379404
rect 91324 379400 91388 379404
rect 91324 379344 91374 379400
rect 91374 379344 91388 379400
rect 91324 379340 91388 379344
rect 92428 379400 92492 379404
rect 92428 379344 92442 379400
rect 92442 379344 92492 379400
rect 92428 379340 92492 379344
rect 93532 379400 93596 379404
rect 93532 379344 93546 379400
rect 93546 379344 93596 379400
rect 93532 379340 93596 379344
rect 96108 379400 96172 379404
rect 96108 379344 96122 379400
rect 96122 379344 96172 379400
rect 96108 379340 96172 379344
rect 98132 379340 98196 379404
rect 98500 379400 98564 379404
rect 98500 379344 98514 379400
rect 98514 379344 98564 379400
rect 98500 379340 98564 379344
rect 101076 379400 101140 379404
rect 101076 379344 101090 379400
rect 101090 379344 101140 379400
rect 101076 379340 101140 379344
rect 103284 379340 103348 379404
rect 105860 379340 105924 379404
rect 108252 379400 108316 379404
rect 108252 379344 108266 379400
rect 108266 379344 108316 379400
rect 108252 379340 108316 379344
rect 108804 379400 108868 379404
rect 108804 379344 108854 379400
rect 108854 379344 108868 379400
rect 108804 379340 108868 379344
rect 111196 379400 111260 379404
rect 111196 379344 111246 379400
rect 111246 379344 111260 379400
rect 111196 379340 111260 379344
rect 112300 379340 112364 379404
rect 113404 379400 113468 379404
rect 113404 379344 113454 379400
rect 113454 379344 113468 379400
rect 113404 379340 113468 379344
rect 114508 379400 114572 379404
rect 114508 379344 114522 379400
rect 114522 379344 114572 379400
rect 114508 379340 114572 379344
rect 117084 379400 117148 379404
rect 117084 379344 117134 379400
rect 117134 379344 117148 379400
rect 117084 379340 117148 379344
rect 141004 379400 141068 379404
rect 141004 379344 141054 379400
rect 141054 379344 141068 379400
rect 141004 379340 141068 379344
rect 148548 379400 148612 379404
rect 148548 379344 148598 379400
rect 148598 379344 148612 379400
rect 148548 379340 148612 379344
rect 150940 379400 151004 379404
rect 150940 379344 150990 379400
rect 150990 379344 151004 379400
rect 150940 379340 151004 379344
rect 153516 379400 153580 379404
rect 153516 379344 153566 379400
rect 153566 379344 153580 379400
rect 153516 379340 153580 379344
rect 183140 379400 183204 379404
rect 183140 379344 183190 379400
rect 183190 379344 183204 379400
rect 183140 379340 183204 379344
rect 199516 379340 199580 379404
rect 246436 379340 246500 379404
rect 247540 379400 247604 379404
rect 247540 379344 247554 379400
rect 247554 379344 247604 379400
rect 247540 379340 247604 379344
rect 248644 379400 248708 379404
rect 248644 379344 248658 379400
rect 248658 379344 248708 379400
rect 248644 379340 248708 379344
rect 250116 379400 250180 379404
rect 250116 379344 250130 379400
rect 250130 379344 250180 379400
rect 250116 379340 250180 379344
rect 251220 379400 251284 379404
rect 251220 379344 251234 379400
rect 251234 379344 251284 379400
rect 251220 379340 251284 379344
rect 252324 379400 252388 379404
rect 252324 379344 252338 379400
rect 252338 379344 252388 379400
rect 252324 379340 252388 379344
rect 253428 379400 253492 379404
rect 253428 379344 253442 379400
rect 253442 379344 253492 379400
rect 253428 379340 253492 379344
rect 257844 379340 257908 379404
rect 261708 379400 261772 379404
rect 261708 379344 261722 379400
rect 261722 379344 261772 379400
rect 261708 379340 261772 379344
rect 268700 379400 268764 379404
rect 268700 379344 268714 379400
rect 268714 379344 268764 379400
rect 268700 379340 268764 379344
rect 271092 379400 271156 379404
rect 271092 379344 271106 379400
rect 271106 379344 271156 379400
rect 271092 379340 271156 379344
rect 272196 379340 272260 379404
rect 273300 379400 273364 379404
rect 273300 379344 273314 379400
rect 273314 379344 273364 379400
rect 273300 379340 273364 379344
rect 274404 379340 274468 379404
rect 275692 379400 275756 379404
rect 275692 379344 275706 379400
rect 275706 379344 275756 379400
rect 275692 379340 275756 379344
rect 276060 379400 276124 379404
rect 276060 379344 276074 379400
rect 276074 379344 276124 379400
rect 276060 379340 276124 379344
rect 276980 379400 277044 379404
rect 276980 379344 276994 379400
rect 276994 379344 277044 379400
rect 276980 379340 277044 379344
rect 278084 379340 278148 379404
rect 285996 379400 286060 379404
rect 285996 379344 286010 379400
rect 286010 379344 286060 379400
rect 285996 379340 286060 379344
rect 288204 379340 288268 379404
rect 290964 379400 291028 379404
rect 290964 379344 290978 379400
rect 290978 379344 291028 379400
rect 290964 379340 291028 379344
rect 293356 379340 293420 379404
rect 295932 379400 295996 379404
rect 295932 379344 295946 379400
rect 295946 379344 295996 379400
rect 295932 379340 295996 379344
rect 298508 379400 298572 379404
rect 298508 379344 298522 379400
rect 298522 379344 298572 379400
rect 298508 379340 298572 379344
rect 300900 379400 300964 379404
rect 300900 379344 300914 379400
rect 300914 379344 300964 379400
rect 300900 379340 300964 379344
rect 303476 379340 303540 379404
rect 305868 379400 305932 379404
rect 305868 379344 305882 379400
rect 305882 379344 305932 379400
rect 305868 379340 305932 379344
rect 311020 379400 311084 379404
rect 311020 379344 311034 379400
rect 311034 379344 311084 379400
rect 311020 379340 311084 379344
rect 313412 379400 313476 379404
rect 313412 379344 313426 379400
rect 313426 379344 313476 379400
rect 313412 379340 313476 379344
rect 315804 379400 315868 379404
rect 315804 379344 315818 379400
rect 315818 379344 315868 379400
rect 315804 379340 315868 379344
rect 318380 379340 318444 379404
rect 323348 379400 323412 379404
rect 323348 379344 323362 379400
rect 323362 379344 323412 379400
rect 323348 379340 323412 379344
rect 325924 379400 325988 379404
rect 325924 379344 325974 379400
rect 325974 379344 325988 379400
rect 325924 379340 325988 379344
rect 343404 379400 343468 379404
rect 343404 379344 343454 379400
rect 343454 379344 343468 379400
rect 343404 379340 343468 379344
rect 396028 379400 396092 379404
rect 396028 379344 396078 379400
rect 396078 379344 396092 379400
rect 396028 379340 396092 379344
rect 397132 379400 397196 379404
rect 397132 379344 397146 379400
rect 397146 379344 397196 379400
rect 397132 379340 397196 379344
rect 404124 379340 404188 379404
rect 406516 379340 406580 379404
rect 407620 379400 407684 379404
rect 407620 379344 407634 379400
rect 407634 379344 407684 379400
rect 407620 379340 407684 379344
rect 408356 379400 408420 379404
rect 408356 379344 408370 379400
rect 408370 379344 408420 379400
rect 408356 379340 408420 379344
rect 411300 379400 411364 379404
rect 411300 379344 411314 379400
rect 411314 379344 411364 379400
rect 411300 379340 411364 379344
rect 412404 379400 412468 379404
rect 412404 379344 412418 379400
rect 412418 379344 412468 379400
rect 412404 379340 412468 379344
rect 413508 379340 413572 379404
rect 414612 379400 414676 379404
rect 414612 379344 414626 379400
rect 414626 379344 414676 379400
rect 414612 379340 414676 379344
rect 423444 379400 423508 379404
rect 423444 379344 423458 379400
rect 423458 379344 423508 379400
rect 423444 379340 423508 379344
rect 426388 379400 426452 379404
rect 426388 379344 426438 379400
rect 426438 379344 426452 379400
rect 426388 379340 426452 379344
rect 427492 379340 427556 379404
rect 435772 379400 435836 379404
rect 435772 379344 435786 379400
rect 435786 379344 435836 379400
rect 435772 379340 435836 379344
rect 439084 379400 439148 379404
rect 439084 379344 439098 379400
rect 439098 379344 439148 379400
rect 439084 379340 439148 379344
rect 448284 379340 448348 379404
rect 451044 379400 451108 379404
rect 451044 379344 451058 379400
rect 451058 379344 451108 379400
rect 451044 379340 451108 379344
rect 453436 379340 453500 379404
rect 455828 379340 455892 379404
rect 458404 379400 458468 379404
rect 458404 379344 458418 379400
rect 458418 379344 458468 379400
rect 458404 379340 458468 379344
rect 460980 379400 461044 379404
rect 460980 379344 460994 379400
rect 460994 379344 461044 379400
rect 460980 379340 461044 379344
rect 463556 379400 463620 379404
rect 463556 379344 463570 379400
rect 463570 379344 463620 379400
rect 463556 379340 463620 379344
rect 475884 379340 475948 379404
rect 78260 379204 78324 379268
rect 80468 379264 80532 379268
rect 80468 379208 80482 379264
rect 80482 379208 80532 379264
rect 80468 379204 80532 379208
rect 81756 379204 81820 379268
rect 95924 379264 95988 379268
rect 95924 379208 95974 379264
rect 95974 379208 95988 379264
rect 79548 379068 79612 379132
rect 95924 379204 95988 379208
rect 99420 379264 99484 379268
rect 99420 379208 99470 379264
rect 99470 379208 99484 379264
rect 99420 379204 99484 379208
rect 102916 379264 102980 379268
rect 102916 379208 102966 379264
rect 102966 379208 102980 379264
rect 102916 379204 102980 379208
rect 105308 379204 105372 379268
rect 109724 379204 109788 379268
rect 278452 379204 278516 379268
rect 279188 379264 279252 379268
rect 279188 379208 279202 379264
rect 279202 379208 279252 379264
rect 279188 379204 279252 379208
rect 280844 379204 280908 379268
rect 283420 379204 283484 379268
rect 398236 379204 398300 379268
rect 403020 379264 403084 379268
rect 403020 379208 403034 379264
rect 403034 379208 403084 379264
rect 403020 379204 403084 379208
rect 405412 379264 405476 379268
rect 405412 379208 405426 379264
rect 405426 379208 405476 379264
rect 405412 379204 405476 379208
rect 410748 379204 410812 379268
rect 415900 379204 415964 379268
rect 416084 379264 416148 379268
rect 416084 379208 416098 379264
rect 416098 379208 416148 379264
rect 416084 379204 416148 379208
rect 437980 379204 438044 379268
rect 473492 379264 473556 379268
rect 473492 379208 473506 379264
rect 473506 379208 473556 379264
rect 473492 379204 473556 379208
rect 480852 379204 480916 379268
rect 503116 379264 503180 379268
rect 503116 379208 503130 379264
rect 503130 379208 503180 379264
rect 503116 379204 503180 379208
rect 503484 379264 503548 379268
rect 503484 379208 503534 379264
rect 503534 379208 503548 379264
rect 503484 379204 503548 379208
rect 78260 378932 78324 378996
rect 239260 379068 239324 379132
rect 399524 379068 399588 379132
rect 44036 378856 44100 378860
rect 44036 378800 44050 378856
rect 44050 378800 44100 378856
rect 44036 378796 44100 378800
rect 83228 378796 83292 378860
rect 241468 378932 241532 378996
rect 376892 378932 376956 378996
rect 433380 379068 433444 379132
rect 465948 379068 466012 379132
rect 478460 378932 478524 378996
rect 483428 378992 483492 378996
rect 483428 378936 483442 378992
rect 483442 378936 483492 378992
rect 483428 378932 483492 378936
rect 94636 378720 94700 378724
rect 94636 378664 94686 378720
rect 94686 378664 94700 378720
rect 94636 378660 94700 378664
rect 97028 378660 97092 378724
rect 138428 378720 138492 378724
rect 138428 378664 138478 378720
rect 138478 378664 138492 378720
rect 138428 378660 138492 378664
rect 241836 378796 241900 378860
rect 248276 378856 248340 378860
rect 248276 378800 248290 378856
rect 248290 378800 248340 378856
rect 248276 378796 248340 378800
rect 402284 378796 402348 378860
rect 468524 378796 468588 378860
rect 470916 378856 470980 378860
rect 470916 378800 470930 378856
rect 470930 378800 470980 378856
rect 470916 378796 470980 378800
rect 238156 378660 238220 378724
rect 400444 378660 400508 378724
rect 418476 378660 418540 378724
rect 426020 378720 426084 378724
rect 426020 378664 426034 378720
rect 426034 378664 426084 378720
rect 426020 378660 426084 378664
rect 428228 378660 428292 378724
rect 115796 378524 115860 378588
rect 240548 378388 240612 378452
rect 241468 378388 241532 378452
rect 241836 378388 241900 378452
rect 253612 378584 253676 378588
rect 253612 378528 253626 378584
rect 253626 378528 253676 378584
rect 253612 378524 253676 378528
rect 258396 378584 258460 378588
rect 258396 378528 258410 378584
rect 258410 378528 258460 378584
rect 258396 378524 258460 378528
rect 260972 378584 261036 378588
rect 260972 378528 260986 378584
rect 260986 378528 261036 378584
rect 260972 378524 261036 378528
rect 263548 378584 263612 378588
rect 263548 378528 263598 378584
rect 263598 378528 263612 378584
rect 263548 378524 263612 378528
rect 265940 378584 266004 378588
rect 265940 378528 265954 378584
rect 265954 378528 266004 378584
rect 265940 378524 266004 378528
rect 268332 378524 268396 378588
rect 273484 378584 273548 378588
rect 273484 378528 273498 378584
rect 273498 378528 273548 378584
rect 273484 378524 273548 378528
rect 320956 378584 321020 378588
rect 320956 378528 320970 378584
rect 320970 378528 321020 378584
rect 320956 378524 321020 378528
rect 417004 378584 417068 378588
rect 417004 378528 417018 378584
rect 417018 378528 417068 378584
rect 417004 378524 417068 378528
rect 436876 378524 436940 378588
rect 343220 378448 343284 378452
rect 343220 378392 343234 378448
rect 343234 378392 343284 378448
rect 343220 378388 343284 378392
rect 104020 378252 104084 378316
rect 107516 378312 107580 378316
rect 107516 378256 107566 378312
rect 107566 378256 107580 378312
rect 107516 378252 107580 378256
rect 118188 378252 118252 378316
rect 244228 378312 244292 378316
rect 244228 378256 244278 378312
rect 244278 378256 244292 378312
rect 244228 378252 244292 378256
rect 250668 378312 250732 378316
rect 250668 378256 250682 378312
rect 250682 378256 250732 378312
rect 250668 378252 250732 378256
rect 262812 378312 262876 378316
rect 262812 378256 262826 378312
rect 262826 378256 262876 378312
rect 262812 378252 262876 378256
rect 266308 378312 266372 378316
rect 266308 378256 266358 378312
rect 266358 378256 266372 378312
rect 266308 378252 266372 378256
rect 267596 378312 267660 378316
rect 267596 378256 267610 378312
rect 267610 378256 267660 378312
rect 267596 378252 267660 378256
rect 431172 378312 431236 378316
rect 431172 378256 431186 378312
rect 431186 378256 431236 378312
rect 431172 378252 431236 378256
rect 84332 378116 84396 378180
rect 100708 378116 100772 378180
rect 101812 378176 101876 378180
rect 101812 378120 101862 378176
rect 101862 378120 101876 378176
rect 101812 378116 101876 378120
rect 106412 378176 106476 378180
rect 106412 378120 106462 378176
rect 106462 378120 106476 378176
rect 106412 378116 106476 378120
rect 183508 378116 183572 378180
rect 211660 378116 211724 378180
rect 308628 378116 308692 378180
rect 199148 377844 199212 377908
rect 217548 377980 217612 378044
rect 376892 378116 376956 378180
rect 410012 378176 410076 378180
rect 410012 378120 410026 378176
rect 410026 378120 410076 378176
rect 410012 378116 410076 378120
rect 418108 378176 418172 378180
rect 418108 378120 418158 378176
rect 418158 378120 418172 378176
rect 418108 378116 418172 378120
rect 420684 378116 420748 378180
rect 421788 378176 421852 378180
rect 421788 378120 421802 378176
rect 421802 378120 421852 378176
rect 421788 378116 421852 378120
rect 423996 378176 424060 378180
rect 423996 378120 424010 378176
rect 424010 378120 424060 378176
rect 423996 378116 424060 378120
rect 425284 378116 425348 378180
rect 428596 378116 428660 378180
rect 429700 378116 429764 378180
rect 432276 378176 432340 378180
rect 432276 378120 432290 378176
rect 432290 378120 432340 378176
rect 432276 378116 432340 378120
rect 359780 377980 359844 378044
rect 216628 377844 216692 377908
rect 213684 376756 213748 376820
rect 370084 376756 370148 376820
rect 377444 376620 377508 376684
rect 209820 375532 209884 375596
rect 213868 375532 213932 375596
rect 57100 375396 57164 375460
rect 208900 375396 208964 375460
rect 210004 375396 210068 375460
rect 214052 375396 214116 375460
rect 377444 375260 377508 375324
rect 375420 375124 375484 375188
rect 217548 374912 217612 374916
rect 217548 374856 217562 374912
rect 217562 374856 217612 374912
rect 217548 374852 217612 374856
rect 377996 374776 378060 374780
rect 377996 374720 378010 374776
rect 378010 374720 378060 374776
rect 377996 374716 378060 374720
rect 199332 371920 199396 371924
rect 199332 371864 199382 371920
rect 199382 371864 199396 371920
rect 199332 371860 199396 371864
rect 178540 358804 178604 358868
rect 179644 358804 179708 358868
rect 190868 358864 190932 358868
rect 190868 358808 190918 358864
rect 190918 358808 190932 358864
rect 190868 358804 190932 358808
rect 338436 358864 338500 358868
rect 338436 358808 338486 358864
rect 338486 358808 338500 358864
rect 338436 358804 338500 358808
rect 339724 358804 339788 358868
rect 350948 358804 351012 358868
rect 498516 358804 498580 358868
rect 499804 358804 499868 358868
rect 510844 358864 510908 358868
rect 510844 358808 510894 358864
rect 510894 358808 510908 358864
rect 510844 358804 510908 358808
rect 54708 282236 54772 282300
rect 95910 273804 95974 273868
rect 113318 273864 113382 273868
rect 113318 273808 113362 273864
rect 113362 273808 113382 273864
rect 113318 273804 113382 273808
rect 274406 273804 274470 273868
rect 133446 273728 133510 273732
rect 133446 273672 133474 273728
rect 133474 273672 133510 273728
rect 133446 273668 133510 273672
rect 135894 273592 135958 273596
rect 135894 273536 135902 273592
rect 135902 273536 135958 273592
rect 135894 273532 135958 273536
rect 138478 273592 138542 273596
rect 138478 273536 138534 273592
rect 138534 273536 138542 273592
rect 138478 273532 138542 273536
rect 140926 273532 140990 273596
rect 143510 273592 143574 273596
rect 143510 273536 143538 273592
rect 143538 273536 143574 273592
rect 143510 273532 143574 273536
rect 145958 273592 146022 273596
rect 145958 273536 145986 273592
rect 145986 273536 146022 273592
rect 145958 273532 146022 273536
rect 266382 273592 266446 273596
rect 266382 273536 266414 273592
rect 266414 273536 266446 273592
rect 266382 273532 266446 273536
rect 269782 273592 269846 273596
rect 269782 273536 269818 273592
rect 269818 273536 269846 273592
rect 269782 273532 269846 273536
rect 271142 273592 271206 273596
rect 271142 273536 271198 273592
rect 271198 273536 271206 273592
rect 271142 273532 271206 273536
rect 283518 273592 283582 273596
rect 283518 273536 283526 273592
rect 283526 273536 283582 273592
rect 283518 273532 283582 273536
rect 421078 273592 421142 273596
rect 421078 273536 421102 273592
rect 421102 273536 421142 273592
rect 421078 273532 421142 273536
rect 422846 273592 422910 273596
rect 422846 273536 422850 273592
rect 422850 273536 422906 273592
rect 422906 273536 422910 273592
rect 422846 273532 422910 273536
rect 427606 273592 427670 273596
rect 427606 273536 427634 273592
rect 427634 273536 427670 273592
rect 427606 273532 427670 273536
rect 445966 273592 446030 273596
rect 445966 273536 445998 273592
rect 445998 273536 446030 273592
rect 445966 273532 446030 273536
rect 273300 273456 273364 273460
rect 273300 273400 273314 273456
rect 273314 273400 273364 273456
rect 273300 273396 273364 273400
rect 377444 273396 377508 273460
rect 377812 273396 377876 273460
rect 378180 273396 378244 273460
rect 215340 273260 215404 273324
rect 217364 273260 217428 273324
rect 250668 273260 250732 273324
rect 359412 273260 359476 273324
rect 430988 273260 431052 273324
rect 76052 273184 76116 273188
rect 76052 273128 76066 273184
rect 76066 273128 76116 273184
rect 76052 273124 76116 273128
rect 77156 273184 77220 273188
rect 77156 273128 77170 273184
rect 77170 273128 77220 273184
rect 77156 273124 77220 273128
rect 90772 273184 90836 273188
rect 90772 273128 90786 273184
rect 90786 273128 90836 273184
rect 90772 273124 90836 273128
rect 93716 273184 93780 273188
rect 93716 273128 93730 273184
rect 93730 273128 93780 273184
rect 93716 273124 93780 273128
rect 101812 273124 101876 273188
rect 198044 273124 198108 273188
rect 318380 273124 318444 273188
rect 359596 273124 359660 273188
rect 483244 273124 483308 273188
rect 47716 272988 47780 273052
rect 97028 272988 97092 273052
rect 196756 272988 196820 273052
rect 298508 273048 298572 273052
rect 298508 272992 298522 273048
rect 298522 272992 298572 273048
rect 94452 272912 94516 272916
rect 94452 272856 94466 272912
rect 94466 272856 94516 272912
rect 94452 272852 94516 272856
rect 95924 272912 95988 272916
rect 95924 272856 95938 272912
rect 95938 272856 95988 272912
rect 95924 272852 95988 272856
rect 98500 272912 98564 272916
rect 98500 272856 98514 272912
rect 98514 272856 98564 272912
rect 98500 272852 98564 272856
rect 285996 272912 286060 272916
rect 285996 272856 286010 272912
rect 286010 272856 286060 272912
rect 285996 272852 286060 272856
rect 288204 272912 288268 272916
rect 288204 272856 288218 272912
rect 288218 272856 288268 272912
rect 288204 272852 288268 272856
rect 290964 272912 291028 272916
rect 290964 272856 290978 272912
rect 290978 272856 291028 272912
rect 290964 272852 291028 272856
rect 293356 272912 293420 272916
rect 293356 272856 293370 272912
rect 293370 272856 293420 272912
rect 293356 272852 293420 272856
rect 295932 272912 295996 272916
rect 295932 272856 295946 272912
rect 295946 272856 295996 272912
rect 295932 272852 295996 272856
rect 298508 272988 298572 272992
rect 377812 272988 377876 273052
rect 423444 273048 423508 273052
rect 423444 272992 423458 273048
rect 423458 272992 423508 273048
rect 305868 272852 305932 272916
rect 423444 272988 423508 272992
rect 425284 273048 425348 273052
rect 425284 272992 425298 273048
rect 425298 272992 425348 273048
rect 425284 272988 425348 272992
rect 426020 273048 426084 273052
rect 426020 272992 426034 273048
rect 426034 272992 426084 273048
rect 426020 272988 426084 272992
rect 428228 273048 428292 273052
rect 428228 272992 428242 273048
rect 428242 272992 428292 273048
rect 428228 272988 428292 272992
rect 468524 273048 468588 273052
rect 468524 272992 468538 273048
rect 468538 272992 468588 273048
rect 468524 272988 468588 272992
rect 423812 272852 423876 272916
rect 470916 272912 470980 272916
rect 470916 272856 470930 272912
rect 470930 272856 470980 272912
rect 470916 272852 470980 272856
rect 478460 272912 478524 272916
rect 478460 272856 478474 272912
rect 478474 272856 478524 272912
rect 478460 272852 478524 272856
rect 103836 272716 103900 272780
rect 300900 272776 300964 272780
rect 300900 272720 300914 272776
rect 300914 272720 300964 272776
rect 300900 272716 300964 272720
rect 303476 272776 303540 272780
rect 303476 272720 303490 272776
rect 303490 272720 303540 272776
rect 303476 272716 303540 272720
rect 473492 272776 473556 272780
rect 473492 272720 473506 272776
rect 473506 272720 473556 272776
rect 473492 272716 473556 272720
rect 480852 272776 480916 272780
rect 480852 272720 480866 272776
rect 480866 272720 480916 272776
rect 480852 272716 480916 272720
rect 118004 272580 118068 272644
rect 311020 272640 311084 272644
rect 311020 272584 311034 272640
rect 311034 272584 311084 272640
rect 311020 272580 311084 272584
rect 320956 272640 321020 272644
rect 320956 272584 320970 272640
rect 320970 272584 321020 272640
rect 320956 272580 321020 272584
rect 475884 272640 475948 272644
rect 475884 272584 475898 272640
rect 475898 272584 475948 272640
rect 475884 272580 475948 272584
rect 486004 272640 486068 272644
rect 486004 272584 486018 272640
rect 486018 272584 486068 272640
rect 486004 272580 486068 272584
rect 108620 272444 108684 272508
rect 83044 272368 83108 272372
rect 83044 272312 83058 272368
rect 83058 272312 83108 272368
rect 83044 272308 83108 272312
rect 100708 272368 100772 272372
rect 100708 272312 100758 272368
rect 100758 272312 100772 272368
rect 100708 272308 100772 272312
rect 99420 272232 99484 272236
rect 99420 272176 99434 272232
rect 99434 272176 99484 272232
rect 99420 272172 99484 272176
rect 265204 272232 265268 272236
rect 265204 272176 265218 272232
rect 265218 272176 265268 272232
rect 265204 272172 265268 272176
rect 401732 272232 401796 272236
rect 401732 272176 401746 272232
rect 401746 272176 401796 272232
rect 401732 272172 401796 272176
rect 415900 272232 415964 272236
rect 415900 272176 415914 272232
rect 415914 272176 415964 272232
rect 415900 272172 415964 272176
rect 416084 272232 416148 272236
rect 416084 272176 416098 272232
rect 416098 272176 416148 272232
rect 416084 272172 416148 272176
rect 455828 272232 455892 272236
rect 455828 272176 455842 272232
rect 455842 272176 455892 272232
rect 455828 272172 455892 272176
rect 51580 271824 51644 271828
rect 51580 271768 51630 271824
rect 51630 271768 51644 271824
rect 51580 271764 51644 271768
rect 53236 271764 53300 271828
rect 83964 271764 84028 271828
rect 98132 271764 98196 271828
rect 102732 271764 102796 271828
rect 105308 271764 105372 271828
rect 107516 271824 107580 271828
rect 107516 271768 107530 271824
rect 107530 271768 107580 271824
rect 107516 271764 107580 271768
rect 114508 271824 114572 271828
rect 114508 271768 114522 271824
rect 114522 271768 114572 271824
rect 114508 271764 114572 271768
rect 123524 271764 123588 271828
rect 125916 271764 125980 271828
rect 130884 271764 130948 271828
rect 150940 271764 151004 271828
rect 154068 271764 154132 271828
rect 158484 271764 158548 271828
rect 263548 271824 263612 271828
rect 263548 271768 263598 271824
rect 263598 271768 263612 271824
rect 263548 271764 263612 271768
rect 270908 271764 270972 271828
rect 272564 271764 272628 271828
rect 276980 271764 277044 271828
rect 278452 271764 278516 271828
rect 280844 271764 280908 271828
rect 308628 271764 308692 271828
rect 343404 271764 343468 271828
rect 428596 271764 428660 271828
rect 431172 271764 431236 271828
rect 432276 271764 432340 271828
rect 433380 271824 433444 271828
rect 433380 271768 433394 271824
rect 433394 271768 433444 271824
rect 433380 271764 433444 271768
rect 435956 271764 436020 271828
rect 438532 271764 438596 271828
rect 443500 271764 443564 271828
rect 448284 271764 448348 271828
rect 451044 271764 451108 271828
rect 453436 271764 453500 271828
rect 458404 271764 458468 271828
rect 81940 271628 82004 271692
rect 101076 271628 101140 271692
rect 111012 271628 111076 271692
rect 120764 271628 120828 271692
rect 128676 271628 128740 271692
rect 155908 271628 155972 271692
rect 160876 271628 160940 271692
rect 163452 271628 163516 271692
rect 166028 271628 166092 271692
rect 183140 271628 183204 271692
rect 315068 271628 315132 271692
rect 465948 271628 466012 271692
rect 503116 271628 503180 271692
rect 79548 271492 79612 271556
rect 115980 271552 116044 271556
rect 115980 271496 115994 271552
rect 115994 271496 116044 271552
rect 115980 271492 116044 271496
rect 118372 271492 118436 271556
rect 217180 271492 217244 271556
rect 273484 271492 273548 271556
rect 276244 271492 276308 271556
rect 460980 271492 461044 271556
rect 78260 271356 78324 271420
rect 103836 271356 103900 271420
rect 113220 271416 113284 271420
rect 113220 271360 113234 271416
rect 113234 271360 113284 271416
rect 113220 271356 113284 271360
rect 236500 271356 236564 271420
rect 260972 271356 261036 271420
rect 268332 271356 268396 271420
rect 343220 271356 343284 271420
rect 377260 271356 377324 271420
rect 408172 271356 408236 271420
rect 433564 271356 433628 271420
rect 440924 271356 440988 271420
rect 105860 271220 105924 271284
rect 108252 271220 108316 271284
rect 119108 271220 119172 271284
rect 258396 271220 258460 271284
rect 265940 271220 266004 271284
rect 275324 271220 275388 271284
rect 278084 271220 278148 271284
rect 396028 271220 396092 271284
rect 439268 271220 439332 271284
rect 503484 271220 503548 271284
rect 112116 271084 112180 271148
rect 248276 271084 248340 271148
rect 253612 271084 253676 271148
rect 256188 271084 256252 271148
rect 313412 271084 313476 271148
rect 397132 271084 397196 271148
rect 410748 271084 410812 271148
rect 413692 271084 413756 271148
rect 418476 271084 418540 271148
rect 80468 270948 80532 271012
rect 88380 271008 88444 271012
rect 88380 270952 88394 271008
rect 88394 270952 88444 271008
rect 88380 270948 88444 270952
rect 90036 270948 90100 271012
rect 115796 270948 115860 271012
rect 325556 270948 325620 271012
rect 462636 270948 462700 271012
rect 86540 270812 86604 270876
rect 88748 270812 88812 270876
rect 93348 270812 93412 270876
rect 106412 270812 106476 270876
rect 116900 270812 116964 270876
rect 148548 270812 148612 270876
rect 254532 270812 254596 270876
rect 279004 270812 279068 270876
rect 406516 270812 406580 270876
rect 434668 270872 434732 270876
rect 434668 270816 434718 270872
rect 434718 270816 434732 270872
rect 434668 270812 434732 270816
rect 436876 270812 436940 270876
rect 438348 270812 438412 270876
rect 244228 270676 244292 270740
rect 251220 270736 251284 270740
rect 251220 270680 251270 270736
rect 251270 270680 251284 270736
rect 251220 270676 251284 270680
rect 255820 270676 255884 270740
rect 260604 270676 260668 270740
rect 411300 270736 411364 270740
rect 411300 270680 411350 270736
rect 411350 270680 411364 270736
rect 411300 270676 411364 270680
rect 429700 270676 429764 270740
rect 435772 270676 435836 270740
rect 84700 270600 84764 270604
rect 84700 270544 84714 270600
rect 84714 270544 84764 270600
rect 84700 270540 84764 270544
rect 87644 270540 87708 270604
rect 91324 270540 91388 270604
rect 109540 270540 109604 270604
rect 111196 270540 111260 270604
rect 183508 270600 183572 270604
rect 183508 270544 183522 270600
rect 183522 270544 183572 270600
rect 183508 270540 183572 270544
rect 237052 270540 237116 270604
rect 238156 270540 238220 270604
rect 242940 270600 243004 270604
rect 242940 270544 242954 270600
rect 242954 270544 243004 270600
rect 242940 270540 243004 270544
rect 245332 270540 245396 270604
rect 246436 270540 246500 270604
rect 247724 270540 247788 270604
rect 248644 270540 248708 270604
rect 250116 270540 250180 270604
rect 252324 270540 252388 270604
rect 253428 270540 253492 270604
rect 256924 270540 256988 270604
rect 258396 270540 258460 270604
rect 259500 270600 259564 270604
rect 259500 270544 259514 270600
rect 259514 270544 259564 270600
rect 259500 270540 259564 270544
rect 262076 270540 262140 270604
rect 262812 270540 262876 270604
rect 263916 270540 263980 270604
rect 267596 270540 267660 270604
rect 268700 270540 268764 270604
rect 397500 270600 397564 270604
rect 397500 270544 397514 270600
rect 397514 270544 397564 270600
rect 397500 270540 397564 270544
rect 399524 270540 399588 270604
rect 400444 270540 400508 270604
rect 403020 270600 403084 270604
rect 403020 270544 403034 270600
rect 403034 270544 403084 270600
rect 403020 270540 403084 270544
rect 404124 270540 404188 270604
rect 405044 270540 405108 270604
rect 407620 270540 407684 270604
rect 408724 270540 408788 270604
rect 410012 270540 410076 270604
rect 412404 270540 412468 270604
rect 413324 270540 413388 270604
rect 414428 270540 414492 270604
rect 417004 270540 417068 270604
rect 418108 270600 418172 270604
rect 418108 270544 418158 270600
rect 418158 270544 418172 270600
rect 418108 270540 418172 270544
rect 420684 270540 420748 270604
rect 421788 270540 421852 270604
rect 57468 270404 57532 270468
rect 91508 270404 91572 270468
rect 323348 270404 323412 270468
rect 241652 270268 241716 270332
rect 419212 270404 419276 270468
rect 240548 270132 240612 270196
rect 217548 269860 217612 269924
rect 239260 269724 239324 269788
rect 426388 269724 426452 269788
rect 44772 269044 44836 269108
rect 44956 268908 45020 268972
rect 217180 268696 217244 268700
rect 217180 268640 217230 268696
rect 217230 268640 217244 268696
rect 217180 268636 217244 268640
rect 377996 264964 378060 265028
rect 54340 253948 54404 254012
rect 339724 253404 339788 253468
rect 179644 253268 179708 253332
rect 499804 253268 499868 253332
rect 178540 253132 178604 253196
rect 190868 253132 190932 253196
rect 350948 253132 351012 253196
rect 338436 252996 338500 253060
rect 498516 252724 498580 252788
rect 510844 252648 510908 252652
rect 510844 252592 510894 252648
rect 510894 252592 510908 252648
rect 510844 252588 510908 252592
rect 377996 252452 378060 252516
rect 53052 201452 53116 201516
rect 57468 175884 57532 175948
rect 57652 175068 57716 175132
rect 57836 166908 57900 166972
rect 202276 166908 202340 166972
rect 356652 166908 356716 166972
rect 47900 166772 47964 166836
rect 93716 166772 93780 166836
rect 96108 166832 96172 166836
rect 96108 166776 96122 166832
rect 96122 166776 96172 166832
rect 96108 166772 96172 166776
rect 98500 166832 98564 166836
rect 98500 166776 98514 166832
rect 98514 166776 98564 166832
rect 98500 166772 98564 166776
rect 101076 166832 101140 166836
rect 101076 166776 101090 166832
rect 101090 166776 101140 166832
rect 101076 166772 101140 166776
rect 105860 166832 105924 166836
rect 105860 166776 105874 166832
rect 105874 166776 105924 166832
rect 105860 166772 105924 166776
rect 108252 166832 108316 166836
rect 108252 166776 108266 166832
rect 108266 166776 108316 166832
rect 108252 166772 108316 166776
rect 138478 166832 138542 166836
rect 138478 166776 138534 166832
rect 138534 166776 138542 166832
rect 138478 166772 138542 166776
rect 140926 166772 140990 166836
rect 143510 166772 143574 166836
rect 145958 166832 146022 166836
rect 145958 166776 145986 166832
rect 145986 166776 146022 166832
rect 145958 166772 146022 166776
rect 202460 166772 202524 166836
rect 305958 166772 306022 166836
rect 313438 166772 313502 166836
rect 418476 166832 418540 166836
rect 418476 166776 418490 166832
rect 418490 166776 418540 166832
rect 418476 166772 418540 166776
rect 421052 166832 421116 166836
rect 421052 166776 421066 166832
rect 421066 166776 421116 166832
rect 421052 166772 421116 166776
rect 428286 166832 428350 166836
rect 428286 166776 428334 166832
rect 428334 166776 428350 166832
rect 428286 166772 428350 166776
rect 431006 166772 431070 166836
rect 433590 166832 433654 166836
rect 433590 166776 433614 166832
rect 433614 166776 433654 166832
rect 433590 166772 433654 166776
rect 470990 166772 471054 166836
rect 473438 166832 473502 166836
rect 473438 166776 473450 166832
rect 473450 166776 473502 166832
rect 473438 166772 473502 166776
rect 475886 166832 475950 166836
rect 475886 166776 475898 166832
rect 475898 166776 475950 166832
rect 475886 166772 475950 166776
rect 478470 166832 478534 166836
rect 478470 166776 478474 166832
rect 478474 166776 478534 166832
rect 478470 166772 478534 166776
rect 480918 166832 480982 166836
rect 480918 166776 480958 166832
rect 480958 166776 480982 166832
rect 480918 166772 480982 166776
rect 163366 166696 163430 166700
rect 163366 166640 163374 166696
rect 163374 166640 163430 166696
rect 163366 166636 163430 166640
rect 203012 166636 203076 166700
rect 288278 166696 288342 166700
rect 288278 166640 288310 166696
rect 288310 166640 288342 166696
rect 288278 166636 288342 166640
rect 290998 166696 291062 166700
rect 290998 166640 291014 166696
rect 291014 166640 291062 166696
rect 290998 166636 291062 166640
rect 483366 166696 483430 166700
rect 483366 166640 483386 166696
rect 483386 166640 483430 166696
rect 483366 166636 483430 166640
rect 485950 166696 486014 166700
rect 485950 166640 485962 166696
rect 485962 166640 486014 166696
rect 485950 166636 486014 166640
rect 111142 166560 111206 166564
rect 111142 166504 111154 166560
rect 111154 166504 111206 166560
rect 111142 166500 111206 166504
rect 116990 166560 117054 166564
rect 116990 166504 117006 166560
rect 117006 166504 117054 166560
rect 116990 166500 117054 166504
rect 148548 166560 148612 166564
rect 148548 166504 148562 166560
rect 148562 166504 148612 166560
rect 148548 166500 148612 166504
rect 213500 166500 213564 166564
rect 303510 166500 303574 166564
rect 434406 166500 434470 166564
rect 503222 166560 503286 166564
rect 503222 166504 503258 166560
rect 503258 166504 503286 166560
rect 503222 166500 503286 166504
rect 153332 166424 153396 166428
rect 153332 166368 153346 166424
rect 153346 166368 153396 166424
rect 153332 166364 153396 166368
rect 196572 166364 196636 166428
rect 260972 166424 261036 166428
rect 260972 166368 260986 166424
rect 260986 166368 261036 166424
rect 260972 166364 261036 166368
rect 265940 166424 266004 166428
rect 265940 166368 265954 166424
rect 265954 166368 266004 166424
rect 265940 166364 266004 166368
rect 293356 166424 293420 166428
rect 293356 166368 293370 166424
rect 293370 166368 293420 166424
rect 270908 166228 270972 166292
rect 285996 166288 286060 166292
rect 293356 166364 293420 166368
rect 298508 166424 298572 166428
rect 298508 166368 298522 166424
rect 298522 166368 298572 166424
rect 298508 166364 298572 166368
rect 285996 166232 286010 166288
rect 286010 166232 286060 166288
rect 285996 166228 286060 166232
rect 295932 166228 295996 166292
rect 423444 166288 423508 166292
rect 423444 166232 423458 166288
rect 423458 166232 423508 166288
rect 423444 166228 423508 166232
rect 81756 165548 81820 165612
rect 85436 165548 85500 165612
rect 92428 165548 92492 165612
rect 95740 165548 95804 165612
rect 99420 165608 99484 165612
rect 99420 165552 99434 165608
rect 99434 165552 99484 165608
rect 99420 165548 99484 165552
rect 103468 165608 103532 165612
rect 103468 165552 103518 165608
rect 103518 165552 103532 165608
rect 103468 165548 103532 165552
rect 109724 165548 109788 165612
rect 111012 165608 111076 165612
rect 111012 165552 111026 165608
rect 111026 165552 111076 165608
rect 111012 165548 111076 165552
rect 113588 165608 113652 165612
rect 113588 165552 113602 165608
rect 113602 165552 113652 165608
rect 113588 165548 113652 165552
rect 115980 165608 116044 165612
rect 115980 165552 115994 165608
rect 115994 165552 116044 165608
rect 115980 165548 116044 165552
rect 118004 165548 118068 165612
rect 118372 165548 118436 165612
rect 120948 165608 121012 165612
rect 120948 165552 120962 165608
rect 120962 165552 121012 165608
rect 120948 165548 121012 165552
rect 123524 165608 123588 165612
rect 123524 165552 123538 165608
rect 123538 165552 123588 165608
rect 123524 165548 123588 165552
rect 125916 165608 125980 165612
rect 125916 165552 125930 165608
rect 125930 165552 125980 165608
rect 125916 165548 125980 165552
rect 128492 165548 128556 165612
rect 130884 165548 130948 165612
rect 133460 165548 133524 165612
rect 135852 165548 135916 165612
rect 150940 165548 151004 165612
rect 183140 165608 183204 165612
rect 183140 165552 183190 165608
rect 183190 165552 183204 165608
rect 183140 165548 183204 165552
rect 183508 165608 183572 165612
rect 183508 165552 183522 165608
rect 183522 165552 183572 165608
rect 183508 165548 183572 165552
rect 218652 165548 218716 165612
rect 236132 165608 236196 165612
rect 236132 165552 236146 165608
rect 236146 165552 236196 165608
rect 236132 165548 236196 165552
rect 239628 165548 239692 165612
rect 243124 165548 243188 165612
rect 247540 165548 247604 165612
rect 256188 165548 256252 165612
rect 258028 165548 258092 165612
rect 261708 165548 261772 165612
rect 278452 165548 278516 165612
rect 280844 165548 280908 165612
rect 283420 165608 283484 165612
rect 283420 165552 283434 165608
rect 283434 165552 283484 165608
rect 283420 165548 283484 165552
rect 300900 165608 300964 165612
rect 300900 165552 300914 165608
rect 300914 165552 300964 165608
rect 300900 165548 300964 165552
rect 308444 165548 308508 165612
rect 320956 165608 321020 165612
rect 320956 165552 320970 165608
rect 320970 165552 321020 165608
rect 320956 165548 321020 165552
rect 325924 165608 325988 165612
rect 325924 165552 325938 165608
rect 325938 165552 325988 165608
rect 325924 165548 325988 165552
rect 343220 165608 343284 165612
rect 343220 165552 343270 165608
rect 343270 165552 343284 165608
rect 343220 165548 343284 165552
rect 343404 165608 343468 165612
rect 343404 165552 343454 165608
rect 343454 165552 343468 165608
rect 343404 165548 343468 165552
rect 398236 165548 398300 165612
rect 401732 165548 401796 165612
rect 405412 165548 405476 165612
rect 408172 165548 408236 165612
rect 415900 165548 415964 165612
rect 416084 165608 416148 165612
rect 416084 165552 416098 165608
rect 416098 165552 416148 165608
rect 416084 165548 416148 165552
rect 419396 165548 419460 165612
rect 423812 165548 423876 165612
rect 427492 165548 427556 165612
rect 429700 165608 429764 165612
rect 429700 165552 429714 165608
rect 429714 165552 429764 165608
rect 429700 165548 429764 165552
rect 435772 165548 435836 165612
rect 435956 165608 436020 165612
rect 435956 165552 435970 165608
rect 435970 165552 436020 165608
rect 435956 165548 436020 165552
rect 437980 165608 438044 165612
rect 437980 165552 437994 165608
rect 437994 165552 438044 165608
rect 437980 165548 438044 165552
rect 438532 165608 438596 165612
rect 438532 165552 438546 165608
rect 438546 165552 438596 165608
rect 438532 165548 438596 165552
rect 439268 165548 439332 165612
rect 440924 165608 440988 165612
rect 440924 165552 440938 165608
rect 440938 165552 440988 165608
rect 440924 165548 440988 165552
rect 443500 165608 443564 165612
rect 443500 165552 443514 165608
rect 443514 165552 443564 165608
rect 443500 165548 443564 165552
rect 445892 165608 445956 165612
rect 445892 165552 445906 165608
rect 445906 165552 445956 165608
rect 445892 165548 445956 165552
rect 448284 165548 448348 165612
rect 451044 165548 451108 165612
rect 453436 165548 453500 165612
rect 455828 165548 455892 165612
rect 458404 165608 458468 165612
rect 458404 165552 458418 165608
rect 458418 165552 458468 165608
rect 458404 165548 458468 165552
rect 503300 165608 503364 165612
rect 503300 165552 503350 165608
rect 503350 165552 503364 165608
rect 503300 165548 503364 165552
rect 158484 165412 158548 165476
rect 166028 165412 166092 165476
rect 198780 165412 198844 165476
rect 205220 165412 205284 165476
rect 315804 165412 315868 165476
rect 468524 165412 468588 165476
rect 155908 165276 155972 165340
rect 206324 165276 206388 165340
rect 311020 165276 311084 165340
rect 465948 165276 466012 165340
rect 160876 165140 160940 165204
rect 208164 165140 208228 165204
rect 263732 165140 263796 165204
rect 265204 165140 265268 165204
rect 268332 165140 268396 165204
rect 272196 165140 272260 165204
rect 275692 165140 275756 165204
rect 276060 165200 276124 165204
rect 276060 165144 276074 165200
rect 276074 165144 276124 165200
rect 276060 165140 276124 165144
rect 279188 165140 279252 165204
rect 374868 165140 374932 165204
rect 463556 165140 463620 165204
rect 119108 165004 119172 165068
rect 273484 165064 273548 165068
rect 273484 165008 273498 165064
rect 273498 165008 273548 165064
rect 273484 165004 273548 165008
rect 379468 165004 379532 165068
rect 426020 165004 426084 165068
rect 432276 165064 432340 165068
rect 432276 165008 432290 165064
rect 432290 165008 432340 165064
rect 432276 165004 432340 165008
rect 114508 164928 114572 164932
rect 114508 164872 114522 164928
rect 114522 164872 114572 164928
rect 114508 164868 114572 164872
rect 248276 164868 248340 164932
rect 250668 164868 250732 164932
rect 253612 164868 253676 164932
rect 258396 164868 258460 164932
rect 413692 164868 413756 164932
rect 436876 164868 436940 164932
rect 88380 164792 88444 164796
rect 88380 164736 88394 164792
rect 88394 164736 88444 164792
rect 88380 164732 88444 164736
rect 90772 164732 90836 164796
rect 200988 164732 201052 164796
rect 323348 164732 323412 164796
rect 410748 164732 410812 164796
rect 112116 164656 112180 164660
rect 112116 164600 112130 164656
rect 112130 164600 112180 164656
rect 112116 164596 112180 164600
rect 115796 164656 115860 164660
rect 115796 164600 115810 164656
rect 115810 164600 115860 164656
rect 115796 164596 115860 164600
rect 460980 164596 461044 164660
rect 97028 164460 97092 164524
rect 113220 164460 113284 164524
rect 421788 164460 421852 164524
rect 431172 164460 431236 164524
rect 77156 164324 77220 164388
rect 101812 164324 101876 164388
rect 103836 164324 103900 164388
rect 244412 164324 244476 164388
rect 252324 164324 252388 164388
rect 260604 164324 260668 164388
rect 266492 164324 266556 164388
rect 274404 164324 274468 164388
rect 397132 164324 397196 164388
rect 404124 164324 404188 164388
rect 412404 164324 412468 164388
rect 76052 164248 76116 164252
rect 76052 164192 76066 164248
rect 76066 164192 76116 164248
rect 76052 164188 76116 164192
rect 78260 164188 78324 164252
rect 79548 164188 79612 164252
rect 80468 164188 80532 164252
rect 83044 164188 83108 164252
rect 84148 164188 84212 164252
rect 86540 164188 86604 164252
rect 87644 164188 87708 164252
rect 88748 164188 88812 164252
rect 90036 164188 90100 164252
rect 91324 164188 91388 164252
rect 93348 164188 93412 164252
rect 94452 164188 94516 164252
rect 98132 164188 98196 164252
rect 100708 164248 100772 164252
rect 100708 164192 100758 164248
rect 100758 164192 100772 164248
rect 100708 164188 100772 164192
rect 102732 164188 102796 164252
rect 105308 164188 105372 164252
rect 106412 164248 106476 164252
rect 106412 164192 106426 164248
rect 106426 164192 106476 164248
rect 106412 164188 106476 164192
rect 107516 164248 107580 164252
rect 107516 164192 107566 164248
rect 107566 164192 107580 164248
rect 107516 164188 107580 164192
rect 108620 164188 108684 164252
rect 237052 164188 237116 164252
rect 238156 164188 238220 164252
rect 240548 164188 240612 164252
rect 241652 164188 241716 164252
rect 245332 164188 245396 164252
rect 246436 164188 246500 164252
rect 248644 164188 248708 164252
rect 250116 164188 250180 164252
rect 251220 164248 251284 164252
rect 251220 164192 251234 164248
rect 251234 164192 251284 164248
rect 251220 164188 251284 164192
rect 253428 164188 253492 164252
rect 254532 164188 254596 164252
rect 255820 164188 255884 164252
rect 256924 164188 256988 164252
rect 259500 164248 259564 164252
rect 259500 164192 259514 164248
rect 259514 164192 259564 164248
rect 259500 164188 259564 164192
rect 262812 164188 262876 164252
rect 263916 164188 263980 164252
rect 267596 164188 267660 164252
rect 268700 164188 268764 164252
rect 269804 164188 269868 164252
rect 271276 164188 271340 164252
rect 273300 164188 273364 164252
rect 276980 164188 277044 164252
rect 278084 164248 278148 164252
rect 278084 164192 278098 164248
rect 278098 164192 278148 164248
rect 278084 164188 278148 164192
rect 57468 164112 57532 164116
rect 57468 164056 57518 164112
rect 57518 164056 57532 164112
rect 57468 164052 57532 164056
rect 214604 164052 214668 164116
rect 318380 164188 318444 164252
rect 396028 164248 396092 164252
rect 396028 164192 396078 164248
rect 396078 164192 396092 164248
rect 396028 164188 396092 164192
rect 399524 164188 399588 164252
rect 400444 164188 400508 164252
rect 403020 164248 403084 164252
rect 403020 164192 403034 164248
rect 403034 164192 403084 164248
rect 403020 164188 403084 164192
rect 406516 164188 406580 164252
rect 407620 164188 407684 164252
rect 408724 164188 408788 164252
rect 410012 164248 410076 164252
rect 410012 164192 410026 164248
rect 410026 164192 410076 164248
rect 410012 164188 410076 164192
rect 411300 164248 411364 164252
rect 411300 164192 411314 164248
rect 411314 164192 411364 164248
rect 411300 164188 411364 164192
rect 413324 164188 413388 164252
rect 414428 164188 414492 164252
rect 417004 164188 417068 164252
rect 418292 164188 418356 164252
rect 420684 164188 420748 164252
rect 422892 164188 422956 164252
rect 425284 164188 425348 164252
rect 426388 164248 426452 164252
rect 426388 164192 426438 164248
rect 426438 164192 426452 164248
rect 426388 164188 426452 164192
rect 428780 164188 428844 164252
rect 433380 164188 433444 164252
rect 207980 163916 208044 163980
rect 217180 162556 217244 162620
rect 360884 149092 360948 149156
rect 217364 148276 217428 148340
rect 377628 148276 377692 148340
rect 57652 147732 57716 147796
rect 377996 146236 378060 146300
rect 379468 146100 379532 146164
rect 377812 145692 377876 145756
rect 379468 145556 379532 145620
rect 510844 145420 510908 145484
rect 178540 144876 178604 144940
rect 179644 144936 179708 144940
rect 179644 144880 179694 144936
rect 179694 144880 179708 144936
rect 179644 144876 179708 144880
rect 190868 144876 190932 144940
rect 338436 144936 338500 144940
rect 338436 144880 338486 144936
rect 338486 144880 338500 144936
rect 338436 144876 338500 144880
rect 339724 144876 339788 144940
rect 350948 144876 351012 144940
rect 498516 144876 498580 144940
rect 499804 144876 499868 144940
rect 57468 140796 57532 140860
rect 46796 67764 46860 67828
rect 214420 68036 214484 68100
rect 376156 68036 376220 68100
rect 219020 60616 219084 60620
rect 219020 60560 219070 60616
rect 219070 60560 219084 60616
rect 219020 60556 219084 60560
rect 77142 59800 77206 59804
rect 77142 59744 77170 59800
rect 77170 59744 77206 59800
rect 77142 59740 77206 59744
rect 83126 59800 83190 59804
rect 83126 59744 83150 59800
rect 83150 59744 83190 59800
rect 83126 59740 83190 59744
rect 101758 59800 101822 59804
rect 101758 59744 101770 59800
rect 101770 59744 101822 59800
rect 101758 59740 101822 59744
rect 103934 59800 103998 59804
rect 103934 59744 103942 59800
rect 103942 59744 103998 59800
rect 103934 59740 103998 59744
rect 107606 59800 107670 59804
rect 107606 59744 107622 59800
rect 107622 59744 107670 59800
rect 107606 59740 107670 59744
rect 113590 59800 113654 59804
rect 113590 59744 113602 59800
rect 113602 59744 113654 59800
rect 113590 59740 113654 59744
rect 236054 59740 236118 59804
rect 237142 59800 237206 59804
rect 237142 59744 237158 59800
rect 237158 59744 237206 59800
rect 237142 59740 237206 59744
rect 255910 59800 255974 59804
rect 255910 59744 255926 59800
rect 255926 59744 255974 59800
rect 255910 59740 255974 59744
rect 256998 59800 257062 59804
rect 256998 59744 257030 59800
rect 257030 59744 257062 59800
rect 256998 59740 257062 59744
rect 262846 59800 262910 59804
rect 262846 59744 262862 59800
rect 262862 59744 262910 59800
rect 262846 59740 262910 59744
rect 396054 59800 396118 59804
rect 396054 59744 396078 59800
rect 396078 59744 396118 59800
rect 396054 59740 396118 59744
rect 397142 59800 397206 59804
rect 397142 59744 397146 59800
rect 397146 59744 397206 59800
rect 397142 59740 397206 59744
rect 403126 59740 403190 59804
rect 416998 59800 417062 59804
rect 416998 59744 417018 59800
rect 417018 59744 417062 59800
rect 416998 59740 417062 59744
rect 422846 59800 422910 59804
rect 422846 59744 422850 59800
rect 422850 59744 422906 59800
rect 422906 59744 422910 59800
rect 422846 59740 422910 59744
rect 423934 59800 423998 59804
rect 423934 59744 423954 59800
rect 423954 59744 423998 59800
rect 423934 59740 423998 59744
rect 94550 59664 94614 59668
rect 94550 59608 94558 59664
rect 94558 59608 94614 59664
rect 94550 59604 94614 59608
rect 96998 59664 97062 59668
rect 96998 59608 97042 59664
rect 97042 59608 97062 59664
rect 96998 59604 97062 59608
rect 98086 59664 98150 59668
rect 98086 59608 98090 59664
rect 98090 59608 98146 59664
rect 98146 59608 98150 59664
rect 98086 59604 98150 59608
rect 100708 59664 100772 59668
rect 100708 59608 100758 59664
rect 100758 59608 100772 59664
rect 100708 59604 100772 59608
rect 102846 59604 102910 59668
rect 95924 59528 95988 59532
rect 95924 59472 95938 59528
rect 95938 59472 95988 59528
rect 95924 59468 95988 59472
rect 46612 59332 46676 59396
rect 105974 59604 106038 59668
rect 108694 59664 108758 59668
rect 108694 59608 108726 59664
rect 108726 59608 108758 59664
rect 108694 59604 108758 59608
rect 260670 59664 260734 59668
rect 260670 59608 260710 59664
rect 260710 59608 260734 59664
rect 260670 59604 260734 59608
rect 308542 59664 308606 59668
rect 308542 59608 308550 59664
rect 308550 59608 308606 59664
rect 308542 59604 308606 59608
rect 315886 59664 315950 59668
rect 315886 59608 315910 59664
rect 315910 59608 315950 59664
rect 315886 59604 315950 59608
rect 404214 59664 404278 59668
rect 404214 59608 404230 59664
rect 404230 59608 404278 59664
rect 404214 59604 404278 59608
rect 413462 59604 413526 59668
rect 423526 59664 423590 59668
rect 423526 59608 423550 59664
rect 423550 59608 423590 59664
rect 423526 59604 423590 59608
rect 111012 59392 111076 59396
rect 111012 59336 111026 59392
rect 111026 59336 111076 59392
rect 111012 59332 111076 59336
rect 200804 59332 200868 59396
rect 263548 59468 263612 59532
rect 259500 59392 259564 59396
rect 259500 59336 259514 59392
rect 259514 59336 259564 59392
rect 259500 59332 259564 59336
rect 261708 59392 261772 59396
rect 261708 59336 261722 59392
rect 261722 59336 261772 59392
rect 261708 59332 261772 59336
rect 410748 59392 410812 59396
rect 410748 59336 410762 59392
rect 410762 59336 410812 59392
rect 410748 59332 410812 59336
rect 414612 59392 414676 59396
rect 414612 59336 414626 59392
rect 414626 59336 414676 59392
rect 414612 59332 414676 59336
rect 416084 59392 416148 59396
rect 416084 59336 416098 59392
rect 416098 59336 416148 59392
rect 416084 59332 416148 59336
rect 418108 59392 418172 59396
rect 418108 59336 418158 59392
rect 418158 59336 418172 59392
rect 418108 59332 418172 59336
rect 419396 59392 419460 59396
rect 419396 59336 419410 59392
rect 419410 59336 419460 59392
rect 419396 59332 419460 59336
rect 420684 59392 420748 59396
rect 420684 59336 420698 59392
rect 420698 59336 420748 59392
rect 420684 59332 420748 59336
rect 421788 59392 421852 59396
rect 421788 59336 421802 59392
rect 421802 59336 421852 59392
rect 421788 59332 421852 59336
rect 428228 59392 428292 59396
rect 428228 59336 428242 59392
rect 428242 59336 428292 59392
rect 428228 59332 428292 59336
rect 54892 59196 54956 59260
rect 143580 59196 143644 59260
rect 148548 59256 148612 59260
rect 148548 59200 148562 59256
rect 148562 59200 148612 59256
rect 148548 59196 148612 59200
rect 150940 59256 151004 59260
rect 150940 59200 150954 59256
rect 150954 59200 151004 59256
rect 150940 59196 151004 59200
rect 198412 59196 198476 59260
rect 276060 59196 276124 59260
rect 279188 59256 279252 59260
rect 279188 59200 279238 59256
rect 279238 59200 279252 59256
rect 279188 59196 279252 59200
rect 290964 59256 291028 59260
rect 290964 59200 290978 59256
rect 290978 59200 291028 59256
rect 290964 59196 291028 59200
rect 300900 59256 300964 59260
rect 300900 59200 300914 59256
rect 300914 59200 300964 59256
rect 300900 59196 300964 59200
rect 320956 59256 321020 59260
rect 320956 59200 320970 59256
rect 320970 59200 321020 59256
rect 320956 59196 321020 59200
rect 325924 59256 325988 59260
rect 325924 59200 325938 59256
rect 325938 59200 325988 59256
rect 325924 59196 325988 59200
rect 357940 59196 358004 59260
rect 480852 59196 480916 59260
rect 53420 59060 53484 59124
rect 140820 59060 140884 59124
rect 206876 59060 206940 59124
rect 280844 59060 280908 59124
rect 373764 59060 373828 59124
rect 483428 59060 483492 59124
rect 52132 58924 52196 58988
rect 138428 58924 138492 58988
rect 212396 58924 212460 58988
rect 285996 58924 286060 58988
rect 371740 58924 371804 58988
rect 473492 58924 473556 58988
rect 475884 58984 475948 58988
rect 475884 58928 475898 58984
rect 475898 58928 475948 58984
rect 475884 58924 475948 58928
rect 55444 58788 55508 58852
rect 135852 58788 135916 58852
rect 198596 58788 198660 58852
rect 268332 58788 268396 58852
rect 364932 58788 364996 58852
rect 453436 58788 453500 58852
rect 468524 58848 468588 58852
rect 468524 58792 468538 58848
rect 468538 58792 468588 58848
rect 468524 58788 468588 58792
rect 59308 58652 59372 58716
rect 120948 58652 121012 58716
rect 197860 58652 197924 58716
rect 253612 58652 253676 58716
rect 374500 58652 374564 58716
rect 463556 58652 463620 58716
rect 48084 58516 48148 58580
rect 108252 58516 108316 58580
rect 200620 58516 200684 58580
rect 250668 58516 250732 58580
rect 375972 58516 376036 58580
rect 458404 58516 458468 58580
rect 59124 58380 59188 58444
rect 101076 58380 101140 58444
rect 217548 58380 217612 58444
rect 257844 58380 257908 58444
rect 85436 58108 85500 58172
rect 92244 58108 92308 58172
rect 99420 58108 99484 58172
rect 128308 58108 128372 58172
rect 153332 58108 153396 58172
rect 265204 58108 265268 58172
rect 272196 58108 272260 58172
rect 275692 58108 275756 58172
rect 398236 58108 398300 58172
rect 401732 58108 401796 58172
rect 405412 58108 405476 58172
rect 455828 58108 455892 58172
rect 83964 57972 84028 58036
rect 76052 57896 76116 57900
rect 76052 57840 76066 57896
rect 76066 57840 76116 57896
rect 76052 57836 76116 57840
rect 78260 57896 78324 57900
rect 78260 57840 78274 57896
rect 78274 57840 78324 57896
rect 78260 57836 78324 57840
rect 79548 57896 79612 57900
rect 79548 57840 79562 57896
rect 79562 57840 79612 57896
rect 79548 57836 79612 57840
rect 80468 57836 80532 57900
rect 81940 57896 82004 57900
rect 81940 57840 81954 57896
rect 81954 57840 82004 57896
rect 81940 57836 82004 57840
rect 86540 57896 86604 57900
rect 86540 57840 86554 57896
rect 86554 57840 86604 57896
rect 86540 57836 86604 57840
rect 87644 57836 87708 57900
rect 88748 57896 88812 57900
rect 88748 57840 88762 57896
rect 88762 57840 88812 57896
rect 88748 57836 88812 57840
rect 90036 57836 90100 57900
rect 90772 57896 90836 57900
rect 90772 57840 90786 57896
rect 90786 57840 90836 57896
rect 90772 57836 90836 57840
rect 91324 57836 91388 57900
rect 93348 57836 93412 57900
rect 93716 57836 93780 57900
rect 109540 57896 109604 57900
rect 109540 57840 109554 57896
rect 109554 57840 109604 57896
rect 109540 57836 109604 57840
rect 112116 57896 112180 57900
rect 112116 57840 112130 57896
rect 112130 57840 112180 57896
rect 112116 57836 112180 57840
rect 114324 57836 114388 57900
rect 115980 57896 116044 57900
rect 115980 57840 115994 57896
rect 115994 57840 116044 57896
rect 115980 57836 116044 57840
rect 116900 57836 116964 57900
rect 123524 57896 123588 57900
rect 123524 57840 123538 57896
rect 123538 57840 123588 57896
rect 123524 57836 123588 57840
rect 125916 57896 125980 57900
rect 125916 57840 125930 57896
rect 125930 57840 125980 57896
rect 125916 57836 125980 57840
rect 130884 57896 130948 57900
rect 130884 57840 130898 57896
rect 130898 57840 130948 57896
rect 130884 57836 130948 57840
rect 133460 57896 133524 57900
rect 133460 57840 133474 57896
rect 133474 57840 133524 57896
rect 133460 57836 133524 57840
rect 145604 57896 145668 57900
rect 145604 57840 145618 57896
rect 145618 57840 145668 57896
rect 145604 57836 145668 57840
rect 183140 57836 183204 57900
rect 238156 57836 238220 57900
rect 239260 57896 239324 57900
rect 239260 57840 239274 57896
rect 239274 57840 239324 57896
rect 239260 57836 239324 57840
rect 240548 57836 240612 57900
rect 241652 57896 241716 57900
rect 241652 57840 241666 57896
rect 241666 57840 241716 57896
rect 241652 57836 241716 57840
rect 242940 57896 243004 57900
rect 242940 57840 242954 57896
rect 242954 57840 243004 57896
rect 242940 57836 243004 57840
rect 244228 57836 244292 57900
rect 245332 57896 245396 57900
rect 245332 57840 245346 57896
rect 245346 57840 245396 57896
rect 245332 57836 245396 57840
rect 246436 57836 246500 57900
rect 247724 57896 247788 57900
rect 247724 57840 247738 57896
rect 247738 57840 247788 57896
rect 247724 57836 247788 57840
rect 248644 57836 248708 57900
rect 250116 57896 250180 57900
rect 250116 57840 250130 57896
rect 250130 57840 250180 57896
rect 250116 57836 250180 57840
rect 256004 57836 256068 57900
rect 57836 57700 57900 57764
rect 118004 57700 118068 57764
rect 183508 57760 183572 57764
rect 183508 57704 183522 57760
rect 183522 57704 183572 57760
rect 183508 57700 183572 57704
rect 205036 57700 205100 57764
rect 258396 57760 258460 57764
rect 258396 57704 258410 57760
rect 258410 57704 258460 57760
rect 258396 57700 258460 57704
rect 263916 57700 263980 57764
rect 270908 57836 270972 57900
rect 271092 57896 271156 57900
rect 271092 57840 271106 57896
rect 271106 57840 271156 57896
rect 271092 57836 271156 57840
rect 273300 57896 273364 57900
rect 273300 57840 273314 57896
rect 273314 57840 273364 57896
rect 273300 57836 273364 57840
rect 276980 57896 277044 57900
rect 276980 57840 276994 57896
rect 276994 57840 277044 57896
rect 276980 57836 277044 57840
rect 288204 57836 288268 57900
rect 293356 57896 293420 57900
rect 293356 57840 293370 57896
rect 293370 57840 293420 57896
rect 293356 57836 293420 57840
rect 295932 57896 295996 57900
rect 295932 57840 295946 57896
rect 295946 57840 295996 57896
rect 295932 57836 295996 57840
rect 298508 57836 298572 57900
rect 303476 57896 303540 57900
rect 303476 57840 303490 57896
rect 303490 57840 303540 57896
rect 303476 57836 303540 57840
rect 305868 57896 305932 57900
rect 305868 57840 305882 57896
rect 305882 57840 305932 57896
rect 305868 57836 305932 57840
rect 311020 57896 311084 57900
rect 311020 57840 311034 57896
rect 311034 57840 311084 57896
rect 311020 57836 311084 57840
rect 313412 57896 313476 57900
rect 313412 57840 313426 57896
rect 313426 57840 313476 57896
rect 313412 57836 313476 57840
rect 318380 57836 318444 57900
rect 323348 57896 323412 57900
rect 323348 57840 323362 57896
rect 323362 57840 323412 57896
rect 323348 57836 323412 57840
rect 343220 57896 343284 57900
rect 343220 57840 343234 57896
rect 343234 57840 343284 57896
rect 343220 57836 343284 57840
rect 343404 57896 343468 57900
rect 343404 57840 343454 57896
rect 343454 57840 343468 57896
rect 343404 57836 343468 57840
rect 399524 57896 399588 57900
rect 399524 57840 399538 57896
rect 399538 57840 399588 57896
rect 399524 57836 399588 57840
rect 400444 57836 400508 57900
rect 406516 57836 406580 57900
rect 407620 57836 407684 57900
rect 408356 57896 408420 57900
rect 408356 57840 408370 57896
rect 408370 57840 408420 57896
rect 408356 57836 408420 57840
rect 408724 57896 408788 57900
rect 408724 57840 408738 57896
rect 408738 57840 408788 57896
rect 408724 57836 408788 57840
rect 410012 57836 410076 57900
rect 412404 57836 412468 57900
rect 415532 57896 415596 57900
rect 415532 57840 415546 57896
rect 415546 57840 415596 57896
rect 415532 57836 415596 57840
rect 425284 57896 425348 57900
rect 425284 57840 425298 57896
rect 425298 57840 425348 57896
rect 425284 57836 425348 57840
rect 426388 57896 426452 57900
rect 426388 57840 426438 57896
rect 426438 57840 426452 57896
rect 426388 57836 426452 57840
rect 428596 57896 428660 57900
rect 428596 57840 428610 57896
rect 428610 57840 428660 57896
rect 428596 57836 428660 57840
rect 429700 57836 429764 57900
rect 431172 57836 431236 57900
rect 432276 57896 432340 57900
rect 432276 57840 432290 57896
rect 432290 57840 432340 57896
rect 432276 57836 432340 57840
rect 433564 57896 433628 57900
rect 433564 57840 433578 57896
rect 433578 57840 433628 57896
rect 433564 57836 433628 57840
rect 434668 57896 434732 57900
rect 434668 57840 434682 57896
rect 434682 57840 434732 57896
rect 434668 57836 434732 57840
rect 435956 57896 436020 57900
rect 435956 57840 435970 57896
rect 435970 57840 436020 57896
rect 435956 57836 436020 57840
rect 436876 57836 436940 57900
rect 438532 57896 438596 57900
rect 438532 57840 438546 57896
rect 438546 57840 438596 57896
rect 438532 57836 438596 57840
rect 445892 57896 445956 57900
rect 445892 57840 445906 57896
rect 445906 57840 445956 57896
rect 445892 57836 445956 57840
rect 460980 57896 461044 57900
rect 460980 57840 460994 57896
rect 460994 57840 461044 57896
rect 267596 57700 267660 57764
rect 268700 57700 268764 57764
rect 269804 57700 269868 57764
rect 274404 57700 274468 57764
rect 358124 57700 358188 57764
rect 443500 57700 443564 57764
rect 57652 57564 57716 57628
rect 58572 57428 58636 57492
rect 106412 57564 106476 57628
rect 111196 57564 111260 57628
rect 113220 57624 113284 57628
rect 113220 57568 113270 57624
rect 113270 57568 113284 57624
rect 113220 57564 113284 57568
rect 115796 57564 115860 57628
rect 119108 57564 119172 57628
rect 155908 57624 155972 57628
rect 155908 57568 155958 57624
rect 155958 57568 155972 57624
rect 155908 57564 155972 57568
rect 160876 57564 160940 57628
rect 165844 57564 165908 57628
rect 213132 57564 213196 57628
rect 278452 57564 278516 57628
rect 374684 57564 374748 57628
rect 460980 57836 461044 57840
rect 465948 57896 466012 57900
rect 465948 57840 465962 57896
rect 465962 57840 466012 57896
rect 465948 57836 466012 57840
rect 470916 57896 470980 57900
rect 470916 57840 470930 57896
rect 470930 57840 470980 57896
rect 470916 57836 470980 57840
rect 478460 57896 478524 57900
rect 478460 57840 478474 57896
rect 478474 57840 478524 57896
rect 478460 57836 478524 57840
rect 486004 57896 486068 57900
rect 486004 57840 486018 57896
rect 486018 57840 486068 57896
rect 486004 57836 486068 57840
rect 503116 57836 503180 57900
rect 503484 57896 503548 57900
rect 503484 57840 503534 57896
rect 503534 57840 503548 57896
rect 503484 57836 503548 57840
rect 105308 57428 105372 57492
rect 203196 57428 203260 57492
rect 251220 57488 251284 57492
rect 251220 57432 251234 57488
rect 251234 57432 251284 57488
rect 251220 57428 251284 57432
rect 252324 57428 252388 57492
rect 253428 57428 253492 57492
rect 254532 57428 254596 57492
rect 266308 57488 266372 57492
rect 266308 57432 266358 57488
rect 266358 57432 266372 57488
rect 266308 57428 266372 57432
rect 370452 57428 370516 57492
rect 433380 57488 433444 57492
rect 433380 57432 433430 57488
rect 433430 57432 433444 57488
rect 433380 57428 433444 57432
rect 435772 57428 435836 57492
rect 438348 57428 438412 57492
rect 58756 57292 58820 57356
rect 98500 57292 98564 57356
rect 213316 57292 213380 57356
rect 265940 57292 266004 57356
rect 379100 57292 379164 57356
rect 448284 57292 448348 57356
rect 50476 57156 50540 57220
rect 88380 57156 88444 57220
rect 103836 57156 103900 57220
rect 202092 57156 202156 57220
rect 248276 57156 248340 57220
rect 378916 57156 378980 57220
rect 418476 57156 418540 57220
rect 427676 57156 427740 57220
rect 430988 57216 431052 57220
rect 430988 57160 431002 57216
rect 431002 57160 431052 57216
rect 430988 57156 431052 57160
rect 440924 57156 440988 57220
rect 58940 57020 59004 57084
rect 96292 57020 96356 57084
rect 215892 57020 215956 57084
rect 260972 57020 261036 57084
rect 378732 57020 378796 57084
rect 413508 57020 413572 57084
rect 411300 56944 411364 56948
rect 411300 56888 411314 56944
rect 411314 56888 411364 56944
rect 411300 56884 411364 56888
rect 55076 56748 55140 56812
rect 118372 56748 118436 56812
rect 163268 56612 163332 56676
rect 216076 56612 216140 56676
rect 283788 56612 283852 56676
rect 360700 56612 360764 56676
rect 451044 56612 451108 56676
rect 53604 56476 53668 56540
rect 219204 56476 219268 56540
rect 426020 56476 426084 56540
rect 50660 56340 50724 56404
rect 158484 56340 158548 56404
rect 219940 56340 220004 56404
rect 421052 56340 421116 56404
rect 55628 56204 55692 56268
rect 201356 56204 201420 56268
rect 273484 56204 273548 56268
rect 377628 56204 377692 56268
rect 439084 56204 439148 56268
rect 217364 56068 217428 56132
rect 277164 56068 277228 56132
rect 379468 56068 379532 56132
rect 377812 55932 377876 55996
rect 48636 55116 48700 55180
rect 50844 54980 50908 55044
rect 52316 54844 52380 54908
rect 57468 54708 57532 54772
rect 204852 3980 204916 4044
rect 210372 3844 210436 3908
rect 363460 3708 363524 3772
rect 367876 3572 367940 3636
rect 363644 3436 363708 3500
rect 367692 3300 367756 3364
rect 206140 3164 206204 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 44955 479636 45021 479637
rect 44955 479572 44956 479636
rect 45020 479572 45021 479636
rect 44955 479571 45021 479572
rect 44771 479500 44837 479501
rect 44771 479436 44772 479500
rect 44836 479436 44837 479500
rect 44771 479435 44837 479436
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 44035 467124 44101 467125
rect 44035 467060 44036 467124
rect 44100 467060 44101 467124
rect 44035 467059 44101 467060
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 44038 378861 44098 467059
rect 44035 378860 44101 378861
rect 44035 378796 44036 378860
rect 44100 378796 44101 378860
rect 44035 378795 44101 378796
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 44774 269109 44834 479435
rect 44771 269108 44837 269109
rect 44771 269044 44772 269108
rect 44836 269044 44837 269108
rect 44771 269043 44837 269044
rect 44958 268973 45018 479571
rect 45234 478894 45854 514338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 633099 60134 636618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 633099 63854 640338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 633099 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 633099 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 633099 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 633099 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 633099 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633099 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 633099 96134 636618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 633099 99854 640338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 633099 103574 644058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 633099 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 633099 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 633099 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 633099 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 54339 632636 54405 632637
rect 54339 632572 54340 632636
rect 54404 632572 54405 632636
rect 54339 632571 54405 632572
rect 53051 632500 53117 632501
rect 53051 632436 53052 632500
rect 53116 632436 53117 632500
rect 53051 632435 53117 632436
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 46795 482900 46861 482901
rect 46795 482836 46796 482900
rect 46860 482836 46861 482900
rect 46795 482835 46861 482836
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 46611 465900 46677 465901
rect 46611 465836 46612 465900
rect 46676 465836 46677 465900
rect 46611 465835 46677 465836
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 44955 268972 45021 268973
rect 44955 268908 44956 268972
rect 45020 268908 45021 268972
rect 44955 268907 45021 268908
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 46614 59397 46674 465835
rect 46798 67829 46858 482835
rect 47715 482764 47781 482765
rect 47715 482700 47716 482764
rect 47780 482700 47781 482764
rect 47715 482699 47781 482700
rect 47718 273053 47778 482699
rect 48954 482614 49574 518058
rect 51947 485484 52013 485485
rect 51947 485420 51948 485484
rect 52012 485420 52013 485484
rect 51947 485419 52013 485420
rect 50291 485212 50357 485213
rect 50291 485148 50292 485212
rect 50356 485148 50357 485212
rect 50291 485147 50357 485148
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 47899 471476 47965 471477
rect 47899 471412 47900 471476
rect 47964 471412 47965 471476
rect 47899 471411 47965 471412
rect 47715 273052 47781 273053
rect 47715 272988 47716 273052
rect 47780 272988 47781 273052
rect 47715 272987 47781 272988
rect 47902 166837 47962 471411
rect 48083 469028 48149 469029
rect 48083 468964 48084 469028
rect 48148 468964 48149 469028
rect 48083 468963 48149 468964
rect 47899 166836 47965 166837
rect 47899 166772 47900 166836
rect 47964 166772 47965 166836
rect 47899 166771 47965 166772
rect 46795 67828 46861 67829
rect 46795 67764 46796 67828
rect 46860 67764 46861 67828
rect 46795 67763 46861 67764
rect 46611 59396 46677 59397
rect 46611 59332 46612 59396
rect 46676 59332 46677 59396
rect 46611 59331 46677 59332
rect 48086 58581 48146 468963
rect 48635 468484 48701 468485
rect 48635 468420 48636 468484
rect 48700 468420 48701 468484
rect 48635 468419 48701 468420
rect 48083 58580 48149 58581
rect 48083 58516 48084 58580
rect 48148 58516 48149 58580
rect 48083 58515 48149 58516
rect 48638 55181 48698 468419
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 50294 379541 50354 485147
rect 50843 468756 50909 468757
rect 50843 468692 50844 468756
rect 50908 468692 50909 468756
rect 50843 468691 50909 468692
rect 50659 468620 50725 468621
rect 50659 468556 50660 468620
rect 50724 468556 50725 468620
rect 50659 468555 50725 468556
rect 50475 466444 50541 466445
rect 50475 466380 50476 466444
rect 50540 466380 50541 466444
rect 50475 466379 50541 466380
rect 50291 379540 50357 379541
rect 50291 379476 50292 379540
rect 50356 379476 50357 379540
rect 50291 379475 50357 379476
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48635 55180 48701 55181
rect 48635 55116 48636 55180
rect 48700 55116 48701 55180
rect 48635 55115 48701 55116
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 50614 49574 86058
rect 50478 57221 50538 466379
rect 50475 57220 50541 57221
rect 50475 57156 50476 57220
rect 50540 57156 50541 57220
rect 50475 57155 50541 57156
rect 50662 56405 50722 468555
rect 50659 56404 50725 56405
rect 50659 56340 50660 56404
rect 50724 56340 50725 56404
rect 50659 56339 50725 56340
rect 50846 55045 50906 468691
rect 51579 465220 51645 465221
rect 51579 465156 51580 465220
rect 51644 465156 51645 465220
rect 51579 465155 51645 465156
rect 51582 271829 51642 465155
rect 51950 388517 52010 485419
rect 52315 468892 52381 468893
rect 52315 468828 52316 468892
rect 52380 468828 52381 468892
rect 52315 468827 52381 468828
rect 52131 465764 52197 465765
rect 52131 465700 52132 465764
rect 52196 465700 52197 465764
rect 52131 465699 52197 465700
rect 51947 388516 52013 388517
rect 51947 388452 51948 388516
rect 52012 388452 52013 388516
rect 51947 388451 52013 388452
rect 51579 271828 51645 271829
rect 51579 271764 51580 271828
rect 51644 271764 51645 271828
rect 51579 271763 51645 271764
rect 52134 58989 52194 465699
rect 52131 58988 52197 58989
rect 52131 58924 52132 58988
rect 52196 58924 52197 58988
rect 52131 58923 52197 58924
rect 50843 55044 50909 55045
rect 50843 54980 50844 55044
rect 50908 54980 50909 55044
rect 50843 54979 50909 54980
rect 52318 54909 52378 468827
rect 53054 201517 53114 632435
rect 53419 485348 53485 485349
rect 53419 485284 53420 485348
rect 53484 485284 53485 485348
rect 53419 485283 53485 485284
rect 53235 484532 53301 484533
rect 53235 484468 53236 484532
rect 53300 484468 53301 484532
rect 53235 484467 53301 484468
rect 53238 271829 53298 484467
rect 53235 271828 53301 271829
rect 53235 271764 53236 271828
rect 53300 271764 53301 271828
rect 53235 271763 53301 271764
rect 53051 201516 53117 201517
rect 53051 201452 53052 201516
rect 53116 201452 53117 201516
rect 53051 201451 53117 201452
rect 53422 59125 53482 485283
rect 53603 484532 53669 484533
rect 53603 484468 53604 484532
rect 53668 484468 53669 484532
rect 53603 484467 53669 484468
rect 53419 59124 53485 59125
rect 53419 59060 53420 59124
rect 53484 59060 53485 59124
rect 53419 59059 53485 59060
rect 53606 56541 53666 484467
rect 54342 254013 54402 632571
rect 55794 597454 56414 632898
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 121683 618492 121749 618493
rect 121683 618428 121684 618492
rect 121748 618428 121749 618492
rect 121683 618427 121749 618428
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 79568 597454 79888 597486
rect 79568 597218 79610 597454
rect 79846 597218 79888 597454
rect 79568 597134 79888 597218
rect 79568 596898 79610 597134
rect 79846 596898 79888 597134
rect 79568 596866 79888 596898
rect 110288 597454 110608 597486
rect 110288 597218 110330 597454
rect 110566 597218 110608 597454
rect 110288 597134 110608 597218
rect 110288 596898 110330 597134
rect 110566 596898 110608 597134
rect 110288 596866 110608 596898
rect 64208 579454 64528 579486
rect 64208 579218 64250 579454
rect 64486 579218 64528 579454
rect 64208 579134 64528 579218
rect 64208 578898 64250 579134
rect 64486 578898 64528 579134
rect 64208 578866 64528 578898
rect 94928 579454 95248 579486
rect 94928 579218 94970 579454
rect 95206 579218 95248 579454
rect 94928 579134 95248 579218
rect 94928 578898 94970 579134
rect 95206 578898 95248 579134
rect 94928 578866 95248 578898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 59514 565174 60134 566000
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 550000 60134 564618
rect 63234 551834 63854 566000
rect 63234 551598 63266 551834
rect 63502 551598 63586 551834
rect 63822 551598 63854 551834
rect 63234 551514 63854 551598
rect 63234 551278 63266 551514
rect 63502 551278 63586 551514
rect 63822 551278 63854 551514
rect 63234 550000 63854 551278
rect 66954 555554 67574 566000
rect 66954 555318 66986 555554
rect 67222 555318 67306 555554
rect 67542 555318 67574 555554
rect 66954 555234 67574 555318
rect 66954 554998 66986 555234
rect 67222 554998 67306 555234
rect 67542 554998 67574 555234
rect 66954 550000 67574 554998
rect 73794 560514 74414 566000
rect 73794 560278 73826 560514
rect 74062 560278 74146 560514
rect 74382 560278 74414 560514
rect 73794 560194 74414 560278
rect 73794 559958 73826 560194
rect 74062 559958 74146 560194
rect 74382 559958 74414 560194
rect 73794 550000 74414 559958
rect 77514 564234 78134 566000
rect 77514 563998 77546 564234
rect 77782 563998 77866 564234
rect 78102 563998 78134 564234
rect 77514 563914 78134 563998
rect 77514 563678 77546 563914
rect 77782 563678 77866 563914
rect 78102 563678 78134 563914
rect 77514 550000 78134 563678
rect 81234 550894 81854 566000
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 550000 81854 550338
rect 84954 554614 85574 566000
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 550000 85574 554058
rect 91794 561454 92414 566000
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 550000 92414 560898
rect 95514 565174 96134 566000
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 550000 96134 564618
rect 99234 551834 99854 566000
rect 99234 551598 99266 551834
rect 99502 551598 99586 551834
rect 99822 551598 99854 551834
rect 99234 551514 99854 551598
rect 99234 551278 99266 551514
rect 99502 551278 99586 551514
rect 99822 551278 99854 551514
rect 99234 550000 99854 551278
rect 102954 555554 103574 566000
rect 102954 555318 102986 555554
rect 103222 555318 103306 555554
rect 103542 555318 103574 555554
rect 102954 555234 103574 555318
rect 102954 554998 102986 555234
rect 103222 554998 103306 555234
rect 103542 554998 103574 555234
rect 102954 550000 103574 554998
rect 109794 560514 110414 566000
rect 109794 560278 109826 560514
rect 110062 560278 110146 560514
rect 110382 560278 110414 560514
rect 109794 560194 110414 560278
rect 109794 559958 109826 560194
rect 110062 559958 110146 560194
rect 110382 559958 110414 560194
rect 109794 550000 110414 559958
rect 113514 564234 114134 566000
rect 113514 563998 113546 564234
rect 113782 563998 113866 564234
rect 114102 563998 114134 564234
rect 113514 563914 114134 563998
rect 113514 563678 113546 563914
rect 113782 563678 113866 563914
rect 114102 563678 114134 563914
rect 113514 550000 114134 563678
rect 117234 550894 117854 566000
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 550000 117854 550338
rect 120954 554614 121574 566000
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 550000 121574 554058
rect 121686 552669 121746 618427
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 121683 552668 121749 552669
rect 121683 552604 121684 552668
rect 121748 552604 121749 552668
rect 121683 552603 121749 552604
rect 127794 550000 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 550000 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 551834 135854 568338
rect 135234 551598 135266 551834
rect 135502 551598 135586 551834
rect 135822 551598 135854 551834
rect 135234 551514 135854 551598
rect 135234 551278 135266 551514
rect 135502 551278 135586 551514
rect 135822 551278 135854 551514
rect 135234 550000 135854 551278
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 555554 139574 572058
rect 138954 555318 138986 555554
rect 139222 555318 139306 555554
rect 139542 555318 139574 555554
rect 138954 555234 139574 555318
rect 138954 554998 138986 555234
rect 139222 554998 139306 555234
rect 139542 554998 139574 555234
rect 138954 550000 139574 554998
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 633099 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 633099 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 633099 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633099 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 633099 168134 636618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 633099 171854 640338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 633099 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 633099 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 633099 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 633099 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 633099 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633099 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 633099 204134 636618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 633099 207854 640338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 633099 211574 644058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 154208 615454 154528 615486
rect 154208 615218 154250 615454
rect 154486 615218 154528 615454
rect 154208 615134 154528 615218
rect 154208 614898 154250 615134
rect 154486 614898 154528 615134
rect 154208 614866 154528 614898
rect 184928 615454 185248 615486
rect 184928 615218 184970 615454
rect 185206 615218 185248 615454
rect 184928 615134 185248 615218
rect 184928 614898 184970 615134
rect 185206 614898 185248 615134
rect 184928 614866 185248 614898
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 169568 597454 169888 597486
rect 169568 597218 169610 597454
rect 169846 597218 169888 597454
rect 169568 597134 169888 597218
rect 169568 596898 169610 597134
rect 169846 596898 169888 597134
rect 169568 596866 169888 596898
rect 200288 597454 200608 597486
rect 200288 597218 200330 597454
rect 200566 597218 200608 597454
rect 200288 597134 200608 597218
rect 200288 596898 200330 597134
rect 200566 596898 200608 597134
rect 200288 596866 200608 596898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 560514 146414 578898
rect 154208 579454 154528 579486
rect 154208 579218 154250 579454
rect 154486 579218 154528 579454
rect 154208 579134 154528 579218
rect 154208 578898 154250 579134
rect 154486 578898 154528 579134
rect 154208 578866 154528 578898
rect 184928 579454 185248 579486
rect 184928 579218 184970 579454
rect 185206 579218 185248 579454
rect 184928 579134 185248 579218
rect 184928 578898 184970 579134
rect 185206 578898 185248 579134
rect 184928 578866 185248 578898
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 145794 560278 145826 560514
rect 146062 560278 146146 560514
rect 146382 560278 146414 560514
rect 145794 560194 146414 560278
rect 145794 559958 145826 560194
rect 146062 559958 146146 560194
rect 146382 559958 146414 560194
rect 145794 550000 146414 559958
rect 149514 564234 150134 566000
rect 149514 563998 149546 564234
rect 149782 563998 149866 564234
rect 150102 563998 150134 564234
rect 149514 563914 150134 563998
rect 149514 563678 149546 563914
rect 149782 563678 149866 563914
rect 150102 563678 150134 563914
rect 149514 550000 150134 563678
rect 153234 550894 153854 566000
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 550000 153854 550338
rect 156954 554614 157574 566000
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 550000 157574 554058
rect 163794 561454 164414 566000
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 550000 164414 560898
rect 167514 565174 168134 566000
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 550000 168134 564618
rect 171234 551834 171854 566000
rect 171234 551598 171266 551834
rect 171502 551598 171586 551834
rect 171822 551598 171854 551834
rect 171234 551514 171854 551598
rect 171234 551278 171266 551514
rect 171502 551278 171586 551514
rect 171822 551278 171854 551514
rect 171234 550000 171854 551278
rect 174954 555554 175574 566000
rect 174954 555318 174986 555554
rect 175222 555318 175306 555554
rect 175542 555318 175574 555554
rect 174954 555234 175574 555318
rect 174954 554998 174986 555234
rect 175222 554998 175306 555234
rect 175542 554998 175574 555234
rect 174954 550000 175574 554998
rect 181794 560514 182414 566000
rect 181794 560278 181826 560514
rect 182062 560278 182146 560514
rect 182382 560278 182414 560514
rect 181794 560194 182414 560278
rect 181794 559958 181826 560194
rect 182062 559958 182146 560194
rect 182382 559958 182414 560194
rect 181794 550000 182414 559958
rect 185514 564234 186134 566000
rect 185514 563998 185546 564234
rect 185782 563998 185866 564234
rect 186102 563998 186134 564234
rect 185514 563914 186134 563998
rect 185514 563678 185546 563914
rect 185782 563678 185866 563914
rect 186102 563678 186134 563914
rect 185514 550000 186134 563678
rect 189234 550894 189854 566000
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 550000 189854 550338
rect 192954 554614 193574 566000
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 550000 193574 554058
rect 199794 561454 200414 566000
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 550000 200414 560898
rect 203514 565174 204134 566000
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 550000 204134 564618
rect 207234 551834 207854 566000
rect 207234 551598 207266 551834
rect 207502 551598 207586 551834
rect 207822 551598 207854 551834
rect 207234 551514 207854 551598
rect 207234 551278 207266 551514
rect 207502 551278 207586 551514
rect 207822 551278 207854 551514
rect 207234 550000 207854 551278
rect 210954 555554 211574 566000
rect 210954 555318 210986 555554
rect 211222 555318 211306 555554
rect 211542 555318 211574 555554
rect 210954 555234 211574 555318
rect 210954 554998 210986 555234
rect 211222 554998 211306 555234
rect 211542 554998 211574 555234
rect 210954 550000 211574 554998
rect 217794 560514 218414 578898
rect 217794 560278 217826 560514
rect 218062 560278 218146 560514
rect 218382 560278 218414 560514
rect 217794 560194 218414 560278
rect 217794 559958 217826 560194
rect 218062 559958 218146 560194
rect 218382 559958 218414 560194
rect 217794 550000 218414 559958
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 564234 222134 582618
rect 221514 563998 221546 564234
rect 221782 563998 221866 564234
rect 222102 563998 222134 564234
rect 221514 563914 222134 563998
rect 221514 563678 221546 563914
rect 221782 563678 221866 563914
rect 222102 563678 222134 563914
rect 221514 550000 222134 563678
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 550000 225854 550338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 550000 229574 554058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 633099 240134 636618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 633099 243854 640338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 633099 247574 644058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 633099 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 633099 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 633099 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 633099 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633099 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 633099 276134 636618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 633099 279854 640338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 633099 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 633099 290414 650898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 633099 294134 654618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 633099 297854 658338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 633099 301574 662058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 235794 597454 236414 632898
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 244208 615454 244528 615486
rect 244208 615218 244250 615454
rect 244486 615218 244528 615454
rect 244208 615134 244528 615218
rect 244208 614898 244250 615134
rect 244486 614898 244528 615134
rect 244208 614866 244528 614898
rect 274928 615454 275248 615486
rect 274928 615218 274970 615454
rect 275206 615218 275248 615454
rect 274928 615134 275248 615218
rect 274928 614898 274970 615134
rect 275206 614898 275248 615134
rect 274928 614866 275248 614898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 259568 597454 259888 597486
rect 259568 597218 259610 597454
rect 259846 597218 259888 597454
rect 259568 597134 259888 597218
rect 259568 596898 259610 597134
rect 259846 596898 259888 597134
rect 259568 596866 259888 596898
rect 290288 597454 290608 597486
rect 290288 597218 290330 597454
rect 290566 597218 290608 597454
rect 290288 597134 290608 597218
rect 290288 596898 290330 597134
rect 290566 596898 290608 597134
rect 290288 596866 290608 596898
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 244208 579454 244528 579486
rect 244208 579218 244250 579454
rect 244486 579218 244528 579454
rect 244208 579134 244528 579218
rect 244208 578898 244250 579134
rect 244486 578898 244528 579134
rect 244208 578866 244528 578898
rect 274928 579454 275248 579486
rect 274928 579218 274970 579454
rect 275206 579218 275248 579454
rect 274928 579134 275248 579218
rect 274928 578898 274970 579134
rect 275206 578898 275248 579134
rect 274928 578866 275248 578898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 550000 236414 560898
rect 239514 565174 240134 566000
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 550000 240134 564618
rect 243234 551834 243854 566000
rect 243234 551598 243266 551834
rect 243502 551598 243586 551834
rect 243822 551598 243854 551834
rect 243234 551514 243854 551598
rect 243234 551278 243266 551514
rect 243502 551278 243586 551514
rect 243822 551278 243854 551514
rect 243234 550000 243854 551278
rect 246954 555554 247574 566000
rect 246954 555318 246986 555554
rect 247222 555318 247306 555554
rect 247542 555318 247574 555554
rect 246954 555234 247574 555318
rect 246954 554998 246986 555234
rect 247222 554998 247306 555234
rect 247542 554998 247574 555234
rect 246954 550000 247574 554998
rect 253794 560514 254414 566000
rect 253794 560278 253826 560514
rect 254062 560278 254146 560514
rect 254382 560278 254414 560514
rect 253794 560194 254414 560278
rect 253794 559958 253826 560194
rect 254062 559958 254146 560194
rect 254382 559958 254414 560194
rect 253794 550000 254414 559958
rect 257514 564234 258134 566000
rect 257514 563998 257546 564234
rect 257782 563998 257866 564234
rect 258102 563998 258134 564234
rect 257514 563914 258134 563998
rect 257514 563678 257546 563914
rect 257782 563678 257866 563914
rect 258102 563678 258134 563914
rect 257514 550000 258134 563678
rect 261234 550894 261854 566000
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 550000 261854 550338
rect 264954 554614 265574 566000
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 550000 265574 554058
rect 271794 561454 272414 566000
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 550000 272414 560898
rect 275514 565174 276134 566000
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 550000 276134 564618
rect 279234 551834 279854 566000
rect 279234 551598 279266 551834
rect 279502 551598 279586 551834
rect 279822 551598 279854 551834
rect 279234 551514 279854 551598
rect 279234 551278 279266 551514
rect 279502 551278 279586 551514
rect 279822 551278 279854 551514
rect 279234 550000 279854 551278
rect 282954 555554 283574 566000
rect 282954 555318 282986 555554
rect 283222 555318 283306 555554
rect 283542 555318 283574 555554
rect 282954 555234 283574 555318
rect 282954 554998 282986 555234
rect 283222 554998 283306 555234
rect 283542 554998 283574 555234
rect 282954 550000 283574 554998
rect 289794 560514 290414 566000
rect 289794 560278 289826 560514
rect 290062 560278 290146 560514
rect 290382 560278 290414 560514
rect 289794 560194 290414 560278
rect 289794 559958 289826 560194
rect 290062 559958 290146 560194
rect 290382 559958 290414 560194
rect 289794 550000 290414 559958
rect 293514 564234 294134 566000
rect 293514 563998 293546 564234
rect 293782 563998 293866 564234
rect 294102 563998 294134 564234
rect 293514 563914 294134 563998
rect 293514 563678 293546 563914
rect 293782 563678 293866 563914
rect 294102 563678 294134 563914
rect 293514 550000 294134 563678
rect 297234 550894 297854 566000
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 550000 297854 550338
rect 300954 554614 301574 566000
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 550000 301574 554058
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 299979 549540 300045 549541
rect 299979 549476 299980 549540
rect 300044 549476 300045 549540
rect 299979 549475 300045 549476
rect 64208 543454 64528 543486
rect 64208 543218 64250 543454
rect 64486 543218 64528 543454
rect 64208 543134 64528 543218
rect 64208 542898 64250 543134
rect 64486 542898 64528 543134
rect 64208 542866 64528 542898
rect 94928 543454 95248 543486
rect 94928 543218 94970 543454
rect 95206 543218 95248 543454
rect 94928 543134 95248 543218
rect 94928 542898 94970 543134
rect 95206 542898 95248 543134
rect 94928 542866 95248 542898
rect 125648 543454 125968 543486
rect 125648 543218 125690 543454
rect 125926 543218 125968 543454
rect 125648 543134 125968 543218
rect 125648 542898 125690 543134
rect 125926 542898 125968 543134
rect 125648 542866 125968 542898
rect 156368 543454 156688 543486
rect 156368 543218 156410 543454
rect 156646 543218 156688 543454
rect 156368 543134 156688 543218
rect 156368 542898 156410 543134
rect 156646 542898 156688 543134
rect 156368 542866 156688 542898
rect 187088 543454 187408 543486
rect 187088 543218 187130 543454
rect 187366 543218 187408 543454
rect 187088 543134 187408 543218
rect 187088 542898 187130 543134
rect 187366 542898 187408 543134
rect 187088 542866 187408 542898
rect 217808 543454 218128 543486
rect 217808 543218 217850 543454
rect 218086 543218 218128 543454
rect 217808 543134 218128 543218
rect 217808 542898 217850 543134
rect 218086 542898 218128 543134
rect 217808 542866 218128 542898
rect 248528 543454 248848 543486
rect 248528 543218 248570 543454
rect 248806 543218 248848 543454
rect 248528 543134 248848 543218
rect 248528 542898 248570 543134
rect 248806 542898 248848 543134
rect 248528 542866 248848 542898
rect 279248 543454 279568 543486
rect 279248 543218 279290 543454
rect 279526 543218 279568 543454
rect 279248 543134 279568 543218
rect 279248 542898 279290 543134
rect 279526 542898 279568 543134
rect 279248 542866 279568 542898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 79568 525454 79888 525486
rect 79568 525218 79610 525454
rect 79846 525218 79888 525454
rect 79568 525134 79888 525218
rect 79568 524898 79610 525134
rect 79846 524898 79888 525134
rect 79568 524866 79888 524898
rect 110288 525454 110608 525486
rect 110288 525218 110330 525454
rect 110566 525218 110608 525454
rect 110288 525134 110608 525218
rect 110288 524898 110330 525134
rect 110566 524898 110608 525134
rect 110288 524866 110608 524898
rect 141008 525454 141328 525486
rect 141008 525218 141050 525454
rect 141286 525218 141328 525454
rect 141008 525134 141328 525218
rect 141008 524898 141050 525134
rect 141286 524898 141328 525134
rect 141008 524866 141328 524898
rect 171728 525454 172048 525486
rect 171728 525218 171770 525454
rect 172006 525218 172048 525454
rect 171728 525134 172048 525218
rect 171728 524898 171770 525134
rect 172006 524898 172048 525134
rect 171728 524866 172048 524898
rect 202448 525454 202768 525486
rect 202448 525218 202490 525454
rect 202726 525218 202768 525454
rect 202448 525134 202768 525218
rect 202448 524898 202490 525134
rect 202726 524898 202768 525134
rect 202448 524866 202768 524898
rect 233168 525454 233488 525486
rect 233168 525218 233210 525454
rect 233446 525218 233488 525454
rect 233168 525134 233488 525218
rect 233168 524898 233210 525134
rect 233446 524898 233488 525134
rect 233168 524866 233488 524898
rect 263888 525454 264208 525486
rect 263888 525218 263930 525454
rect 264166 525218 264208 525454
rect 263888 525134 264208 525218
rect 263888 524898 263930 525134
rect 264166 524898 264208 525134
rect 263888 524866 264208 524898
rect 294608 525454 294928 525486
rect 294608 525218 294650 525454
rect 294886 525218 294928 525454
rect 294608 525134 294928 525218
rect 294608 524898 294650 525134
rect 294886 524898 294928 525134
rect 294608 524866 294928 524898
rect 299982 522613 300042 549475
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 299979 522612 300045 522613
rect 299979 522548 299980 522612
rect 300044 522548 300045 522612
rect 299979 522547 300045 522548
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 54707 485620 54773 485621
rect 54707 485556 54708 485620
rect 54772 485556 54773 485620
rect 54707 485555 54773 485556
rect 54710 282301 54770 485555
rect 55075 466308 55141 466309
rect 55075 466244 55076 466308
rect 55140 466244 55141 466308
rect 55075 466243 55141 466244
rect 54891 466036 54957 466037
rect 54891 465972 54892 466036
rect 54956 465972 54957 466036
rect 54891 465971 54957 465972
rect 54707 282300 54773 282301
rect 54707 282236 54708 282300
rect 54772 282236 54773 282300
rect 54707 282235 54773 282236
rect 54339 254012 54405 254013
rect 54339 253948 54340 254012
rect 54404 253948 54405 254012
rect 54339 253947 54405 253948
rect 54894 59261 54954 465971
rect 54891 59260 54957 59261
rect 54891 59196 54892 59260
rect 54956 59196 54957 59260
rect 54891 59195 54957 59196
rect 55078 56813 55138 466243
rect 55443 466172 55509 466173
rect 55443 466108 55444 466172
rect 55508 466108 55509 466172
rect 55443 466107 55509 466108
rect 55446 58853 55506 466107
rect 55627 465220 55693 465221
rect 55627 465156 55628 465220
rect 55692 465156 55693 465220
rect 55627 465155 55693 465156
rect 55443 58852 55509 58853
rect 55443 58788 55444 58852
rect 55508 58788 55509 58852
rect 55443 58787 55509 58788
rect 55075 56812 55141 56813
rect 55075 56748 55076 56812
rect 55140 56748 55141 56812
rect 55075 56747 55141 56748
rect 53603 56540 53669 56541
rect 53603 56476 53604 56540
rect 53668 56476 53669 56540
rect 53603 56475 53669 56476
rect 55630 56269 55690 465155
rect 55794 453454 56414 488898
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 206139 486436 206205 486437
rect 206139 486372 206140 486436
rect 206204 486372 206205 486436
rect 206139 486371 206205 486372
rect 59307 485756 59373 485757
rect 59307 485692 59308 485756
rect 59372 485692 59373 485756
rect 59307 485691 59373 485692
rect 57835 485076 57901 485077
rect 57835 485012 57836 485076
rect 57900 485012 57901 485076
rect 57835 485011 57901 485012
rect 57467 479908 57533 479909
rect 57467 479844 57468 479908
rect 57532 479844 57533 479908
rect 57467 479843 57533 479844
rect 57099 479772 57165 479773
rect 57099 479708 57100 479772
rect 57164 479708 57165 479772
rect 57099 479707 57165 479708
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 57102 375461 57162 479707
rect 57099 375460 57165 375461
rect 57099 375396 57100 375460
rect 57164 375396 57165 375460
rect 57099 375395 57165 375396
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57470 270469 57530 479843
rect 57651 388516 57717 388517
rect 57651 388452 57652 388516
rect 57716 388452 57717 388516
rect 57651 388451 57717 388452
rect 57467 270468 57533 270469
rect 57467 270404 57468 270468
rect 57532 270404 57533 270468
rect 57467 270403 57533 270404
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 57467 175948 57533 175949
rect 57467 175884 57468 175948
rect 57532 175884 57533 175948
rect 57467 175883 57533 175884
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57470 164117 57530 175883
rect 57654 175133 57714 388451
rect 57651 175132 57717 175133
rect 57651 175068 57652 175132
rect 57716 175068 57717 175132
rect 57651 175067 57717 175068
rect 57838 166973 57898 485011
rect 59123 484940 59189 484941
rect 59123 484876 59124 484940
rect 59188 484876 59189 484940
rect 59123 484875 59189 484876
rect 58939 469844 59005 469845
rect 58939 469780 58940 469844
rect 59004 469780 59005 469844
rect 58939 469779 59005 469780
rect 58755 469164 58821 469165
rect 58755 469100 58756 469164
rect 58820 469100 58821 469164
rect 58755 469099 58821 469100
rect 58571 465628 58637 465629
rect 58571 465564 58572 465628
rect 58636 465564 58637 465628
rect 58571 465563 58637 465564
rect 57835 166972 57901 166973
rect 57835 166908 57836 166972
rect 57900 166908 57901 166972
rect 57835 166907 57901 166908
rect 57467 164116 57533 164117
rect 57467 164052 57468 164116
rect 57532 164052 57533 164116
rect 57467 164051 57533 164052
rect 57470 161490 57530 164051
rect 57470 161430 57898 161490
rect 57651 147796 57717 147797
rect 57651 147732 57652 147796
rect 57716 147732 57717 147796
rect 57651 147731 57717 147732
rect 57467 140860 57533 140861
rect 57467 140796 57468 140860
rect 57532 140796 57533 140860
rect 57467 140795 57533 140796
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55627 56268 55693 56269
rect 55627 56204 55628 56268
rect 55692 56204 55693 56268
rect 55627 56203 55693 56204
rect 52315 54908 52381 54909
rect 52315 54844 52316 54908
rect 52380 54844 52381 54908
rect 52315 54843 52381 54844
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 56898
rect 57470 54773 57530 140795
rect 57654 57629 57714 147731
rect 57838 57765 57898 161430
rect 57835 57764 57901 57765
rect 57835 57700 57836 57764
rect 57900 57700 57901 57764
rect 57835 57699 57901 57700
rect 57651 57628 57717 57629
rect 57651 57564 57652 57628
rect 57716 57564 57717 57628
rect 57651 57563 57717 57564
rect 58574 57493 58634 465563
rect 58571 57492 58637 57493
rect 58571 57428 58572 57492
rect 58636 57428 58637 57492
rect 58571 57427 58637 57428
rect 58758 57357 58818 469099
rect 58755 57356 58821 57357
rect 58755 57292 58756 57356
rect 58820 57292 58821 57356
rect 58755 57291 58821 57292
rect 58942 57085 59002 469779
rect 59126 58445 59186 484875
rect 59310 58717 59370 485691
rect 59514 476114 60134 486000
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 60134 476114
rect 59514 475794 60134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 60134 475794
rect 59514 466308 60134 475558
rect 63234 477954 63854 486000
rect 63234 477718 63266 477954
rect 63502 477718 63586 477954
rect 63822 477718 63854 477954
rect 63234 477634 63854 477718
rect 63234 477398 63266 477634
rect 63502 477398 63586 477634
rect 63822 477398 63854 477634
rect 60227 467260 60293 467261
rect 60227 467196 60228 467260
rect 60292 467196 60293 467260
rect 60227 467195 60293 467196
rect 60230 464810 60290 467195
rect 63234 466308 63854 477398
rect 66954 481674 67574 486000
rect 66954 481438 66986 481674
rect 67222 481438 67306 481674
rect 67542 481438 67574 481674
rect 66954 481354 67574 481438
rect 66954 481118 66986 481354
rect 67222 481118 67306 481354
rect 67542 481118 67574 481354
rect 66954 466308 67574 481118
rect 73794 471454 74414 486000
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 466308 74414 470898
rect 77514 475174 78134 486000
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 466308 78134 474618
rect 81234 478894 81854 486000
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 466308 81854 478338
rect 84954 482614 85574 486000
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 466308 85574 482058
rect 91794 472394 92414 486000
rect 91794 472158 91826 472394
rect 92062 472158 92146 472394
rect 92382 472158 92414 472394
rect 91794 472074 92414 472158
rect 91794 471838 91826 472074
rect 92062 471838 92146 472074
rect 92382 471838 92414 472074
rect 91794 466308 92414 471838
rect 95514 476114 96134 486000
rect 95514 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 96134 476114
rect 95514 475794 96134 475878
rect 95514 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 96134 475794
rect 95514 466308 96134 475558
rect 99234 477954 99854 486000
rect 99234 477718 99266 477954
rect 99502 477718 99586 477954
rect 99822 477718 99854 477954
rect 99234 477634 99854 477718
rect 99234 477398 99266 477634
rect 99502 477398 99586 477634
rect 99822 477398 99854 477634
rect 99234 466308 99854 477398
rect 102954 481674 103574 486000
rect 102954 481438 102986 481674
rect 103222 481438 103306 481674
rect 103542 481438 103574 481674
rect 102954 481354 103574 481438
rect 102954 481118 102986 481354
rect 103222 481118 103306 481354
rect 103542 481118 103574 481354
rect 102954 466308 103574 481118
rect 109794 471454 110414 486000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 466308 110414 470898
rect 113514 475174 114134 486000
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 466308 114134 474618
rect 117234 478894 117854 486000
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 466308 117854 478338
rect 120954 482614 121574 486000
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 466308 121574 482058
rect 127794 472394 128414 486000
rect 127794 472158 127826 472394
rect 128062 472158 128146 472394
rect 128382 472158 128414 472394
rect 127794 472074 128414 472158
rect 127794 471838 127826 472074
rect 128062 471838 128146 472074
rect 128382 471838 128414 472074
rect 127794 466308 128414 471838
rect 131514 476114 132134 486000
rect 131514 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 132134 476114
rect 131514 475794 132134 475878
rect 131514 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 132134 475794
rect 131514 466308 132134 475558
rect 135234 477954 135854 486000
rect 135234 477718 135266 477954
rect 135502 477718 135586 477954
rect 135822 477718 135854 477954
rect 135234 477634 135854 477718
rect 135234 477398 135266 477634
rect 135502 477398 135586 477634
rect 135822 477398 135854 477634
rect 135234 466308 135854 477398
rect 138954 481674 139574 486000
rect 138954 481438 138986 481674
rect 139222 481438 139306 481674
rect 139542 481438 139574 481674
rect 138954 481354 139574 481438
rect 138954 481118 138986 481354
rect 139222 481118 139306 481354
rect 139542 481118 139574 481354
rect 138954 466308 139574 481118
rect 145794 471454 146414 486000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 466308 146414 470898
rect 149514 475174 150134 486000
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 466308 150134 474618
rect 153234 478894 153854 486000
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 466308 153854 478338
rect 156954 482614 157574 486000
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 466308 157574 482058
rect 163794 472394 164414 486000
rect 163794 472158 163826 472394
rect 164062 472158 164146 472394
rect 164382 472158 164414 472394
rect 163794 472074 164414 472158
rect 163794 471838 163826 472074
rect 164062 471838 164146 472074
rect 164382 471838 164414 472074
rect 163794 466308 164414 471838
rect 167514 476114 168134 486000
rect 167514 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 168134 476114
rect 167514 475794 168134 475878
rect 167514 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 168134 475794
rect 167514 466308 168134 475558
rect 171234 477954 171854 486000
rect 171234 477718 171266 477954
rect 171502 477718 171586 477954
rect 171822 477718 171854 477954
rect 171234 477634 171854 477718
rect 171234 477398 171266 477634
rect 171502 477398 171586 477634
rect 171822 477398 171854 477634
rect 171234 466308 171854 477398
rect 174954 481674 175574 486000
rect 174954 481438 174986 481674
rect 175222 481438 175306 481674
rect 175542 481438 175574 481674
rect 174954 481354 175574 481438
rect 174954 481118 174986 481354
rect 175222 481118 175306 481354
rect 175542 481118 175574 481354
rect 174954 466308 175574 481118
rect 181794 471454 182414 486000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 179643 467260 179709 467261
rect 179643 467196 179644 467260
rect 179708 467196 179709 467260
rect 179643 467195 179709 467196
rect 178355 466580 178421 466581
rect 178355 466516 178356 466580
rect 178420 466516 178421 466580
rect 178355 466515 178421 466516
rect 59862 464750 60290 464810
rect 178358 464810 178418 466515
rect 179646 464810 179706 467195
rect 181794 466308 182414 470898
rect 185514 475174 186134 486000
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 466308 186134 474618
rect 189234 478894 189854 486000
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 466308 189854 478338
rect 192954 482614 193574 486000
rect 196755 485756 196821 485757
rect 196755 485692 196756 485756
rect 196820 485692 196821 485756
rect 196755 485691 196821 485692
rect 196571 485484 196637 485485
rect 196571 485420 196572 485484
rect 196636 485420 196637 485484
rect 196571 485419 196637 485420
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 190867 466580 190933 466581
rect 190867 466516 190868 466580
rect 190932 466516 190933 466580
rect 190867 466515 190933 466516
rect 190870 464810 190930 466515
rect 192954 466308 193574 482058
rect 178358 464750 178524 464810
rect 179646 464750 179748 464810
rect 59862 381037 59922 464750
rect 178464 464202 178524 464750
rect 179688 464202 179748 464750
rect 190840 464750 190930 464810
rect 190840 464202 190900 464750
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 60952 399454 61300 399486
rect 60952 399218 61008 399454
rect 61244 399218 61300 399454
rect 60952 399134 61300 399218
rect 60952 398898 61008 399134
rect 61244 398898 61300 399134
rect 60952 398866 61300 398898
rect 195320 399454 195668 399486
rect 195320 399218 195376 399454
rect 195612 399218 195668 399454
rect 195320 399134 195668 399218
rect 195320 398898 195376 399134
rect 195612 398898 195668 399134
rect 195320 398866 195668 398898
rect 59859 381036 59925 381037
rect 59859 380972 59860 381036
rect 59924 380972 59925 381036
rect 59859 380971 59925 380972
rect 76056 380493 76116 381106
rect 77144 380629 77204 381106
rect 77141 380628 77207 380629
rect 77141 380564 77142 380628
rect 77206 380564 77207 380628
rect 77141 380563 77207 380564
rect 76051 380492 76117 380493
rect 76051 380428 76052 380492
rect 76116 380428 76117 380492
rect 78232 380490 78292 381106
rect 79592 380490 79652 381106
rect 80544 380490 80604 381106
rect 81768 380490 81828 381106
rect 78232 380430 78322 380490
rect 76051 380427 76117 380428
rect 78262 379269 78322 380430
rect 79550 380430 79652 380490
rect 80470 380430 80604 380490
rect 81758 380430 81828 380490
rect 83128 380490 83188 381106
rect 84216 380490 84276 381106
rect 85440 380490 85500 381106
rect 83128 380430 83290 380490
rect 84216 380430 84394 380490
rect 79550 379405 79610 380430
rect 79547 379404 79613 379405
rect 79547 379340 79548 379404
rect 79612 379340 79613 379404
rect 79547 379339 79613 379340
rect 78259 379268 78325 379269
rect 78259 379204 78260 379268
rect 78324 379204 78325 379268
rect 78259 379203 78325 379204
rect 59514 368114 60134 379000
rect 59514 367878 59546 368114
rect 59782 367878 59866 368114
rect 60102 367878 60134 368114
rect 59514 367794 60134 367878
rect 59514 367558 59546 367794
rect 59782 367558 59866 367794
rect 60102 367558 60134 367794
rect 59514 359308 60134 367558
rect 63234 369954 63854 379000
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 63854 369954
rect 63234 369634 63854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 63854 369634
rect 63234 359308 63854 369398
rect 66954 373674 67574 379000
rect 66954 373438 66986 373674
rect 67222 373438 67306 373674
rect 67542 373438 67574 373674
rect 66954 373354 67574 373438
rect 66954 373118 66986 373354
rect 67222 373118 67306 373354
rect 67542 373118 67574 373354
rect 66954 359308 67574 373118
rect 73794 363454 74414 379000
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 359308 74414 362898
rect 77514 367174 78134 379000
rect 78262 378997 78322 379203
rect 79550 379133 79610 379339
rect 80470 379269 80530 380430
rect 81758 379269 81818 380430
rect 80467 379268 80533 379269
rect 80467 379204 80468 379268
rect 80532 379204 80533 379268
rect 80467 379203 80533 379204
rect 81755 379268 81821 379269
rect 81755 379204 81756 379268
rect 81820 379204 81821 379268
rect 81755 379203 81821 379204
rect 79547 379132 79613 379133
rect 79547 379068 79548 379132
rect 79612 379068 79613 379132
rect 79547 379067 79613 379068
rect 78259 378996 78325 378997
rect 78259 378932 78260 378996
rect 78324 378932 78325 378996
rect 78259 378931 78325 378932
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 359308 78134 366618
rect 81234 370894 81854 379000
rect 83230 378861 83290 380430
rect 83227 378860 83293 378861
rect 83227 378796 83228 378860
rect 83292 378796 83293 378860
rect 83227 378795 83293 378796
rect 84334 378181 84394 380430
rect 85438 380430 85500 380490
rect 86528 380490 86588 381106
rect 87616 380490 87676 381106
rect 88296 380490 88356 381106
rect 88704 380490 88764 381106
rect 90064 380490 90124 381106
rect 86528 380430 86602 380490
rect 87616 380430 87706 380490
rect 88296 380430 88442 380490
rect 88704 380430 88810 380490
rect 85438 379405 85498 380430
rect 86542 379405 86602 380430
rect 87646 379405 87706 380430
rect 88382 379405 88442 380430
rect 88750 379405 88810 380430
rect 90038 380430 90124 380490
rect 90744 380490 90804 381106
rect 91288 380490 91348 381106
rect 92376 380490 92436 381106
rect 93464 380901 93524 381106
rect 93461 380900 93527 380901
rect 93461 380836 93462 380900
rect 93526 380836 93527 380900
rect 93461 380835 93527 380836
rect 93600 380490 93660 381106
rect 90744 380430 90834 380490
rect 91288 380430 91386 380490
rect 92376 380430 92490 380490
rect 90038 379405 90098 380430
rect 90774 379405 90834 380430
rect 91326 379405 91386 380430
rect 92430 379405 92490 380430
rect 93534 380430 93660 380490
rect 94552 380490 94612 381106
rect 95912 380490 95972 381106
rect 96048 380490 96108 381106
rect 97000 380490 97060 381106
rect 98088 380490 98148 381106
rect 98496 380490 98556 381106
rect 99448 380490 99508 381106
rect 94552 380430 94698 380490
rect 95912 380430 95986 380490
rect 96048 380430 96170 380490
rect 97000 380430 97090 380490
rect 98088 380430 98194 380490
rect 98496 380430 98562 380490
rect 93534 379405 93594 380430
rect 85435 379404 85501 379405
rect 85435 379340 85436 379404
rect 85500 379340 85501 379404
rect 85435 379339 85501 379340
rect 86539 379404 86605 379405
rect 86539 379340 86540 379404
rect 86604 379340 86605 379404
rect 86539 379339 86605 379340
rect 87643 379404 87709 379405
rect 87643 379340 87644 379404
rect 87708 379340 87709 379404
rect 87643 379339 87709 379340
rect 88379 379404 88445 379405
rect 88379 379340 88380 379404
rect 88444 379340 88445 379404
rect 88379 379339 88445 379340
rect 88747 379404 88813 379405
rect 88747 379340 88748 379404
rect 88812 379340 88813 379404
rect 88747 379339 88813 379340
rect 90035 379404 90101 379405
rect 90035 379340 90036 379404
rect 90100 379340 90101 379404
rect 90035 379339 90101 379340
rect 90771 379404 90837 379405
rect 90771 379340 90772 379404
rect 90836 379340 90837 379404
rect 90771 379339 90837 379340
rect 91323 379404 91389 379405
rect 91323 379340 91324 379404
rect 91388 379340 91389 379404
rect 91323 379339 91389 379340
rect 92427 379404 92493 379405
rect 92427 379340 92428 379404
rect 92492 379340 92493 379404
rect 92427 379339 92493 379340
rect 93531 379404 93597 379405
rect 93531 379340 93532 379404
rect 93596 379340 93597 379404
rect 93531 379339 93597 379340
rect 84331 378180 84397 378181
rect 84331 378116 84332 378180
rect 84396 378116 84397 378180
rect 84331 378115 84397 378116
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 359308 81854 370338
rect 84954 374614 85574 379000
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 359308 85574 374058
rect 91794 364394 92414 379000
rect 94638 378725 94698 380430
rect 95926 379269 95986 380430
rect 96110 379405 96170 380430
rect 96107 379404 96173 379405
rect 96107 379340 96108 379404
rect 96172 379340 96173 379404
rect 96107 379339 96173 379340
rect 95923 379268 95989 379269
rect 95923 379204 95924 379268
rect 95988 379204 95989 379268
rect 95923 379203 95989 379204
rect 94635 378724 94701 378725
rect 94635 378660 94636 378724
rect 94700 378660 94701 378724
rect 94635 378659 94701 378660
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 92414 364394
rect 91794 364074 92414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 92414 364074
rect 91794 359308 92414 363838
rect 95514 368114 96134 379000
rect 97030 378725 97090 380430
rect 98134 379405 98194 380430
rect 98502 379405 98562 380430
rect 99422 380430 99508 380490
rect 100672 380490 100732 381106
rect 101080 380490 101140 381106
rect 100672 380430 100770 380490
rect 98131 379404 98197 379405
rect 98131 379340 98132 379404
rect 98196 379340 98197 379404
rect 98131 379339 98197 379340
rect 98499 379404 98565 379405
rect 98499 379340 98500 379404
rect 98564 379340 98565 379404
rect 98499 379339 98565 379340
rect 99422 379269 99482 380430
rect 99419 379268 99485 379269
rect 99419 379204 99420 379268
rect 99484 379204 99485 379268
rect 99419 379203 99485 379204
rect 97027 378724 97093 378725
rect 97027 378660 97028 378724
rect 97092 378660 97093 378724
rect 97027 378659 97093 378660
rect 95514 367878 95546 368114
rect 95782 367878 95866 368114
rect 96102 367878 96134 368114
rect 95514 367794 96134 367878
rect 95514 367558 95546 367794
rect 95782 367558 95866 367794
rect 96102 367558 96134 367794
rect 95514 359308 96134 367558
rect 99234 369954 99854 379000
rect 100710 378181 100770 380430
rect 101078 380430 101140 380490
rect 101760 380490 101820 381106
rect 102848 380490 102908 381106
rect 103528 380490 103588 381106
rect 101760 380430 101874 380490
rect 102848 380430 102978 380490
rect 101078 379405 101138 380430
rect 101075 379404 101141 379405
rect 101075 379340 101076 379404
rect 101140 379340 101141 379404
rect 101075 379339 101141 379340
rect 101814 378181 101874 380430
rect 102918 379269 102978 380430
rect 103286 380430 103588 380490
rect 103936 380490 103996 381106
rect 105296 380490 105356 381106
rect 105976 380490 106036 381106
rect 103936 380430 104082 380490
rect 105296 380430 105370 380490
rect 103286 379405 103346 380430
rect 103283 379404 103349 379405
rect 103283 379340 103284 379404
rect 103348 379340 103349 379404
rect 103283 379339 103349 379340
rect 102915 379268 102981 379269
rect 102915 379204 102916 379268
rect 102980 379204 102981 379268
rect 102915 379203 102981 379204
rect 100707 378180 100773 378181
rect 100707 378116 100708 378180
rect 100772 378116 100773 378180
rect 100707 378115 100773 378116
rect 101811 378180 101877 378181
rect 101811 378116 101812 378180
rect 101876 378116 101877 378180
rect 101811 378115 101877 378116
rect 99234 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 99854 369954
rect 99234 369634 99854 369718
rect 99234 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 99854 369634
rect 99234 359308 99854 369398
rect 102954 373674 103574 379000
rect 104022 378317 104082 380430
rect 105310 379269 105370 380430
rect 105862 380430 106036 380490
rect 106384 380490 106444 381106
rect 107608 380490 107668 381106
rect 108288 380490 108348 381106
rect 106384 380430 106474 380490
rect 105862 379405 105922 380430
rect 105859 379404 105925 379405
rect 105859 379340 105860 379404
rect 105924 379340 105925 379404
rect 105859 379339 105925 379340
rect 105307 379268 105373 379269
rect 105307 379204 105308 379268
rect 105372 379204 105373 379268
rect 105307 379203 105373 379204
rect 104019 378316 104085 378317
rect 104019 378252 104020 378316
rect 104084 378252 104085 378316
rect 104019 378251 104085 378252
rect 106414 378181 106474 380430
rect 107518 380430 107668 380490
rect 108254 380430 108348 380490
rect 108696 380490 108756 381106
rect 109784 380490 109844 381106
rect 111008 380901 111068 381106
rect 111005 380900 111071 380901
rect 111005 380836 111006 380900
rect 111070 380836 111071 380900
rect 111005 380835 111071 380836
rect 108696 380430 108866 380490
rect 107518 378317 107578 380430
rect 108254 379405 108314 380430
rect 108806 379405 108866 380430
rect 109726 380430 109844 380490
rect 111144 380490 111204 381106
rect 112232 380490 112292 381106
rect 113320 380490 113380 381106
rect 113592 380901 113652 381106
rect 113589 380900 113655 380901
rect 113589 380836 113590 380900
rect 113654 380836 113655 380900
rect 113589 380835 113655 380836
rect 114408 380490 114468 381106
rect 115768 380490 115828 381106
rect 116040 380901 116100 381106
rect 116037 380900 116103 380901
rect 116037 380836 116038 380900
rect 116102 380836 116103 380900
rect 116037 380835 116103 380836
rect 116992 380490 117052 381106
rect 118080 380490 118140 381106
rect 118488 380901 118548 381106
rect 118485 380900 118551 380901
rect 118485 380836 118486 380900
rect 118550 380836 118551 380900
rect 118485 380835 118551 380836
rect 119168 380490 119228 381106
rect 120936 380901 120996 381106
rect 123520 380901 123580 381106
rect 125968 380901 126028 381106
rect 120933 380900 120999 380901
rect 120933 380836 120934 380900
rect 120998 380836 120999 380900
rect 120933 380835 120999 380836
rect 123517 380900 123583 380901
rect 123517 380836 123518 380900
rect 123582 380836 123583 380900
rect 123517 380835 123583 380836
rect 125965 380900 126031 380901
rect 125965 380836 125966 380900
rect 126030 380836 126031 380900
rect 125965 380835 126031 380836
rect 111144 380430 111258 380490
rect 112232 380430 112362 380490
rect 113320 380430 113466 380490
rect 114408 380430 114570 380490
rect 115768 380430 115858 380490
rect 116992 380430 117146 380490
rect 118080 380430 118250 380490
rect 108251 379404 108317 379405
rect 108251 379340 108252 379404
rect 108316 379340 108317 379404
rect 108251 379339 108317 379340
rect 108803 379404 108869 379405
rect 108803 379340 108804 379404
rect 108868 379340 108869 379404
rect 108803 379339 108869 379340
rect 109726 379269 109786 380430
rect 111198 379405 111258 380430
rect 112302 379405 112362 380430
rect 113406 379405 113466 380430
rect 114510 379405 114570 380430
rect 111195 379404 111261 379405
rect 111195 379340 111196 379404
rect 111260 379340 111261 379404
rect 111195 379339 111261 379340
rect 112299 379404 112365 379405
rect 112299 379340 112300 379404
rect 112364 379340 112365 379404
rect 112299 379339 112365 379340
rect 113403 379404 113469 379405
rect 113403 379340 113404 379404
rect 113468 379340 113469 379404
rect 113403 379339 113469 379340
rect 114507 379404 114573 379405
rect 114507 379340 114508 379404
rect 114572 379340 114573 379404
rect 114507 379339 114573 379340
rect 109723 379268 109789 379269
rect 109723 379204 109724 379268
rect 109788 379204 109789 379268
rect 109723 379203 109789 379204
rect 107515 378316 107581 378317
rect 107515 378252 107516 378316
rect 107580 378252 107581 378316
rect 107515 378251 107581 378252
rect 106411 378180 106477 378181
rect 106411 378116 106412 378180
rect 106476 378116 106477 378180
rect 106411 378115 106477 378116
rect 102954 373438 102986 373674
rect 103222 373438 103306 373674
rect 103542 373438 103574 373674
rect 102954 373354 103574 373438
rect 102954 373118 102986 373354
rect 103222 373118 103306 373354
rect 103542 373118 103574 373354
rect 102954 359308 103574 373118
rect 109794 363454 110414 379000
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 359308 110414 362898
rect 113514 367174 114134 379000
rect 115798 378589 115858 380430
rect 117086 379405 117146 380430
rect 117083 379404 117149 379405
rect 117083 379340 117084 379404
rect 117148 379340 117149 379404
rect 117083 379339 117149 379340
rect 115795 378588 115861 378589
rect 115795 378524 115796 378588
rect 115860 378524 115861 378588
rect 115795 378523 115861 378524
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 359308 114134 366618
rect 117234 370894 117854 379000
rect 118190 378317 118250 380430
rect 119110 380430 119228 380490
rect 128280 380490 128340 381106
rect 131000 380901 131060 381106
rect 133448 380901 133508 381106
rect 135896 380901 135956 381106
rect 130997 380900 131063 380901
rect 130997 380836 130998 380900
rect 131062 380836 131063 380900
rect 130997 380835 131063 380836
rect 133445 380900 133511 380901
rect 133445 380836 133446 380900
rect 133510 380836 133511 380900
rect 133445 380835 133511 380836
rect 135893 380900 135959 380901
rect 135893 380836 135894 380900
rect 135958 380836 135959 380900
rect 135893 380835 135959 380836
rect 138480 380490 138540 381106
rect 128280 380430 128370 380490
rect 119110 380221 119170 380430
rect 128310 380357 128370 380430
rect 138430 380430 138540 380490
rect 140928 380490 140988 381106
rect 143512 380901 143572 381106
rect 145960 380901 146020 381106
rect 143509 380900 143575 380901
rect 143509 380836 143510 380900
rect 143574 380836 143575 380900
rect 143509 380835 143575 380836
rect 145957 380900 146023 380901
rect 145957 380836 145958 380900
rect 146022 380836 146023 380900
rect 145957 380835 146023 380836
rect 148544 380490 148604 381106
rect 150992 380490 151052 381106
rect 140928 380430 141066 380490
rect 148544 380430 148610 380490
rect 128307 380356 128373 380357
rect 128307 380292 128308 380356
rect 128372 380292 128373 380356
rect 128307 380291 128373 380292
rect 119107 380220 119173 380221
rect 119107 380156 119108 380220
rect 119172 380156 119173 380220
rect 119107 380155 119173 380156
rect 118187 378316 118253 378317
rect 118187 378252 118188 378316
rect 118252 378252 118253 378316
rect 118187 378251 118253 378252
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 359308 117854 370338
rect 120954 374614 121574 379000
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 359308 121574 374058
rect 127794 364394 128414 379000
rect 127794 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 128414 364394
rect 127794 364074 128414 364158
rect 127794 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 128414 364074
rect 127794 359308 128414 363838
rect 131514 368114 132134 379000
rect 131514 367878 131546 368114
rect 131782 367878 131866 368114
rect 132102 367878 132134 368114
rect 131514 367794 132134 367878
rect 131514 367558 131546 367794
rect 131782 367558 131866 367794
rect 132102 367558 132134 367794
rect 131514 359308 132134 367558
rect 135234 369954 135854 379000
rect 138430 378725 138490 380430
rect 141006 379405 141066 380430
rect 148550 379405 148610 380430
rect 150942 380430 151052 380490
rect 153440 380490 153500 381106
rect 155888 380490 155948 381106
rect 158472 380901 158532 381106
rect 160920 380901 160980 381106
rect 163368 380901 163428 381106
rect 165952 380901 166012 381106
rect 158469 380900 158535 380901
rect 158469 380836 158470 380900
rect 158534 380836 158535 380900
rect 158469 380835 158535 380836
rect 160917 380900 160983 380901
rect 160917 380836 160918 380900
rect 160982 380836 160983 380900
rect 160917 380835 160983 380836
rect 163365 380900 163431 380901
rect 163365 380836 163366 380900
rect 163430 380836 163431 380900
rect 163365 380835 163431 380836
rect 165949 380900 166015 380901
rect 165949 380836 165950 380900
rect 166014 380836 166015 380900
rect 165949 380835 166015 380836
rect 183224 380490 183284 381106
rect 153440 380430 153578 380490
rect 155888 380430 155970 380490
rect 150942 379405 151002 380430
rect 153518 379405 153578 380430
rect 155910 380357 155970 380430
rect 183142 380430 183284 380490
rect 183360 380490 183420 381106
rect 183360 380430 183570 380490
rect 155907 380356 155973 380357
rect 155907 380292 155908 380356
rect 155972 380292 155973 380356
rect 155907 380291 155973 380292
rect 183142 379405 183202 380430
rect 141003 379404 141069 379405
rect 141003 379340 141004 379404
rect 141068 379340 141069 379404
rect 141003 379339 141069 379340
rect 148547 379404 148613 379405
rect 148547 379340 148548 379404
rect 148612 379340 148613 379404
rect 148547 379339 148613 379340
rect 150939 379404 151005 379405
rect 150939 379340 150940 379404
rect 151004 379340 151005 379404
rect 150939 379339 151005 379340
rect 153515 379404 153581 379405
rect 153515 379340 153516 379404
rect 153580 379340 153581 379404
rect 153515 379339 153581 379340
rect 183139 379404 183205 379405
rect 183139 379340 183140 379404
rect 183204 379340 183205 379404
rect 183139 379339 183205 379340
rect 138427 378724 138493 378725
rect 138427 378660 138428 378724
rect 138492 378660 138493 378724
rect 138427 378659 138493 378660
rect 135234 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 135854 369954
rect 135234 369634 135854 369718
rect 135234 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 135854 369634
rect 135234 359308 135854 369398
rect 138954 373674 139574 379000
rect 138954 373438 138986 373674
rect 139222 373438 139306 373674
rect 139542 373438 139574 373674
rect 138954 373354 139574 373438
rect 138954 373118 138986 373354
rect 139222 373118 139306 373354
rect 139542 373118 139574 373354
rect 138954 359308 139574 373118
rect 145794 363454 146414 379000
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 359308 146414 362898
rect 149514 367174 150134 379000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 359308 150134 366618
rect 153234 370894 153854 379000
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 359308 153854 370338
rect 156954 374614 157574 379000
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 359308 157574 374058
rect 163794 364394 164414 379000
rect 163794 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 164414 364394
rect 163794 364074 164414 364158
rect 163794 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 164414 364074
rect 163794 359308 164414 363838
rect 167514 368114 168134 379000
rect 167514 367878 167546 368114
rect 167782 367878 167866 368114
rect 168102 367878 168134 368114
rect 167514 367794 168134 367878
rect 167514 367558 167546 367794
rect 167782 367558 167866 367794
rect 168102 367558 168134 367794
rect 167514 359308 168134 367558
rect 171234 369954 171854 379000
rect 171234 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 171854 369954
rect 171234 369634 171854 369718
rect 171234 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 171854 369634
rect 171234 359308 171854 369398
rect 174954 373674 175574 379000
rect 174954 373438 174986 373674
rect 175222 373438 175306 373674
rect 175542 373438 175574 373674
rect 174954 373354 175574 373438
rect 174954 373118 174986 373354
rect 175222 373118 175306 373354
rect 175542 373118 175574 373354
rect 174954 359308 175574 373118
rect 181794 363454 182414 379000
rect 183510 378181 183570 380430
rect 183507 378180 183573 378181
rect 183507 378116 183508 378180
rect 183572 378116 183573 378180
rect 183507 378115 183573 378116
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 359308 182414 362898
rect 185514 367174 186134 379000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 359308 186134 366618
rect 189234 370894 189854 379000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 359308 189854 370338
rect 192954 374614 193574 379000
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 359308 193574 374058
rect 178539 358868 178605 358869
rect 178539 358804 178540 358868
rect 178604 358804 178605 358868
rect 178539 358803 178605 358804
rect 179643 358868 179709 358869
rect 179643 358804 179644 358868
rect 179708 358804 179709 358868
rect 179643 358803 179709 358804
rect 190867 358868 190933 358869
rect 190867 358804 190868 358868
rect 190932 358804 190933 358868
rect 190867 358803 190933 358804
rect 178542 358050 178602 358803
rect 178464 357990 178602 358050
rect 179646 358050 179706 358803
rect 190870 358050 190930 358803
rect 179646 357990 179748 358050
rect 178464 357202 178524 357990
rect 179688 357202 179748 357990
rect 190840 357990 190930 358050
rect 190840 357202 190900 357990
rect 60272 345454 60620 345486
rect 60272 345218 60328 345454
rect 60564 345218 60620 345454
rect 60272 345134 60620 345218
rect 60272 344898 60328 345134
rect 60564 344898 60620 345134
rect 60272 344866 60620 344898
rect 196000 345454 196348 345486
rect 196000 345218 196056 345454
rect 196292 345218 196348 345454
rect 196000 345134 196348 345218
rect 196000 344898 196056 345134
rect 196292 344898 196348 345134
rect 196000 344866 196348 344898
rect 60952 327454 61300 327486
rect 60952 327218 61008 327454
rect 61244 327218 61300 327454
rect 60952 327134 61300 327218
rect 60952 326898 61008 327134
rect 61244 326898 61300 327134
rect 60952 326866 61300 326898
rect 195320 327454 195668 327486
rect 195320 327218 195376 327454
rect 195612 327218 195668 327454
rect 195320 327134 195668 327218
rect 195320 326898 195376 327134
rect 195612 326898 195668 327134
rect 195320 326866 195668 326898
rect 60272 309454 60620 309486
rect 60272 309218 60328 309454
rect 60564 309218 60620 309454
rect 60272 309134 60620 309218
rect 60272 308898 60328 309134
rect 60564 308898 60620 309134
rect 60272 308866 60620 308898
rect 196000 309454 196348 309486
rect 196000 309218 196056 309454
rect 196292 309218 196348 309454
rect 196000 309134 196348 309218
rect 196000 308898 196056 309134
rect 196292 308898 196348 309134
rect 196000 308866 196348 308898
rect 60952 291454 61300 291486
rect 60952 291218 61008 291454
rect 61244 291218 61300 291454
rect 60952 291134 61300 291218
rect 60952 290898 61008 291134
rect 61244 290898 61300 291134
rect 60952 290866 61300 290898
rect 195320 291454 195668 291486
rect 195320 291218 195376 291454
rect 195612 291218 195668 291454
rect 195320 291134 195668 291218
rect 195320 290898 195376 291134
rect 195612 290898 195668 291134
rect 195320 290866 195668 290898
rect 76056 273730 76116 274040
rect 76054 273670 76116 273730
rect 77144 273730 77204 274040
rect 78232 273730 78292 274040
rect 79592 273730 79652 274040
rect 80544 273730 80604 274040
rect 77144 273670 77218 273730
rect 78232 273670 78322 273730
rect 76054 273189 76114 273670
rect 77158 273189 77218 273670
rect 76051 273188 76117 273189
rect 76051 273124 76052 273188
rect 76116 273124 76117 273188
rect 76051 273123 76117 273124
rect 77155 273188 77221 273189
rect 77155 273124 77156 273188
rect 77220 273124 77221 273188
rect 77155 273123 77221 273124
rect 59514 260114 60134 272000
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 60134 260114
rect 59514 259794 60134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 60134 259794
rect 59514 252308 60134 259558
rect 63234 261954 63854 272000
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 63854 261954
rect 63234 261634 63854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 63854 261634
rect 63234 252308 63854 261398
rect 66954 265674 67574 272000
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 67574 265674
rect 66954 265354 67574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 67574 265354
rect 66954 252308 67574 265118
rect 73794 255454 74414 272000
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 252308 74414 254898
rect 77514 259174 78134 272000
rect 78262 271421 78322 273670
rect 79550 273670 79652 273730
rect 80470 273670 80604 273730
rect 81768 273730 81828 274040
rect 83128 273730 83188 274040
rect 84216 273730 84276 274040
rect 85440 273730 85500 274040
rect 81768 273670 82002 273730
rect 79550 271557 79610 273670
rect 79547 271556 79613 271557
rect 79547 271492 79548 271556
rect 79612 271492 79613 271556
rect 79547 271491 79613 271492
rect 78259 271420 78325 271421
rect 78259 271356 78260 271420
rect 78324 271356 78325 271420
rect 78259 271355 78325 271356
rect 80470 271013 80530 273670
rect 80467 271012 80533 271013
rect 80467 270948 80468 271012
rect 80532 270948 80533 271012
rect 80467 270947 80533 270948
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 252308 78134 258618
rect 81234 262894 81854 272000
rect 81942 271693 82002 273670
rect 83046 273670 83188 273730
rect 83966 273670 84276 273730
rect 84702 273670 85500 273730
rect 86528 273730 86588 274040
rect 87616 273730 87676 274040
rect 88296 273730 88356 274040
rect 88704 273730 88764 274040
rect 90064 273730 90124 274040
rect 86528 273670 86602 273730
rect 87616 273670 87706 273730
rect 88296 273670 88442 273730
rect 88704 273670 88810 273730
rect 83046 272373 83106 273670
rect 83043 272372 83109 272373
rect 83043 272308 83044 272372
rect 83108 272308 83109 272372
rect 83043 272307 83109 272308
rect 83966 271829 84026 273670
rect 83963 271828 84029 271829
rect 83963 271764 83964 271828
rect 84028 271764 84029 271828
rect 83963 271763 84029 271764
rect 81939 271692 82005 271693
rect 81939 271628 81940 271692
rect 82004 271628 82005 271692
rect 81939 271627 82005 271628
rect 84702 270605 84762 273670
rect 84699 270604 84765 270605
rect 84699 270540 84700 270604
rect 84764 270540 84765 270604
rect 84699 270539 84765 270540
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 252308 81854 262338
rect 84954 266614 85574 272000
rect 86542 270877 86602 273670
rect 86539 270876 86605 270877
rect 86539 270812 86540 270876
rect 86604 270812 86605 270876
rect 86539 270811 86605 270812
rect 87646 270605 87706 273670
rect 88382 271013 88442 273670
rect 88379 271012 88445 271013
rect 88379 270948 88380 271012
rect 88444 270948 88445 271012
rect 88379 270947 88445 270948
rect 88750 270877 88810 273670
rect 90038 273670 90124 273730
rect 90744 273730 90804 274040
rect 91288 273730 91348 274040
rect 92376 273730 92436 274040
rect 93464 273730 93524 274040
rect 90744 273670 90834 273730
rect 91288 273670 91386 273730
rect 90038 271013 90098 273670
rect 90774 273189 90834 273670
rect 90771 273188 90837 273189
rect 90771 273124 90772 273188
rect 90836 273124 90837 273188
rect 90771 273123 90837 273124
rect 90035 271012 90101 271013
rect 90035 270948 90036 271012
rect 90100 270948 90101 271012
rect 90035 270947 90101 270948
rect 88747 270876 88813 270877
rect 88747 270812 88748 270876
rect 88812 270812 88813 270876
rect 88747 270811 88813 270812
rect 91326 270605 91386 273670
rect 91510 273670 92436 273730
rect 93350 273670 93524 273730
rect 93600 273730 93660 274040
rect 94552 273730 94612 274040
rect 95912 273869 95972 274040
rect 95909 273868 95975 273869
rect 95909 273804 95910 273868
rect 95974 273804 95975 273868
rect 95909 273803 95975 273804
rect 96048 273730 96108 274040
rect 93600 273670 93778 273730
rect 87643 270604 87709 270605
rect 87643 270540 87644 270604
rect 87708 270540 87709 270604
rect 87643 270539 87709 270540
rect 91323 270604 91389 270605
rect 91323 270540 91324 270604
rect 91388 270540 91389 270604
rect 91323 270539 91389 270540
rect 91510 270469 91570 273670
rect 91507 270468 91573 270469
rect 91507 270404 91508 270468
rect 91572 270404 91573 270468
rect 91507 270403 91573 270404
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 252308 85574 266058
rect 91794 256394 92414 272000
rect 93350 270877 93410 273670
rect 93718 273189 93778 273670
rect 94454 273670 94612 273730
rect 95926 273670 96108 273730
rect 97000 273730 97060 274040
rect 98088 273730 98148 274040
rect 98496 273730 98556 274040
rect 99448 273730 99508 274040
rect 97000 273670 97090 273730
rect 98088 273670 98194 273730
rect 98496 273670 98562 273730
rect 93715 273188 93781 273189
rect 93715 273124 93716 273188
rect 93780 273124 93781 273188
rect 93715 273123 93781 273124
rect 94454 272917 94514 273670
rect 95926 272917 95986 273670
rect 97030 273053 97090 273670
rect 97027 273052 97093 273053
rect 97027 272988 97028 273052
rect 97092 272988 97093 273052
rect 97027 272987 97093 272988
rect 94451 272916 94517 272917
rect 94451 272852 94452 272916
rect 94516 272852 94517 272916
rect 94451 272851 94517 272852
rect 95923 272916 95989 272917
rect 95923 272852 95924 272916
rect 95988 272852 95989 272916
rect 95923 272851 95989 272852
rect 93347 270876 93413 270877
rect 93347 270812 93348 270876
rect 93412 270812 93413 270876
rect 93347 270811 93413 270812
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 92414 256394
rect 91794 256074 92414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 92414 256074
rect 91794 252308 92414 255838
rect 95514 260114 96134 272000
rect 98134 271829 98194 273670
rect 98502 272917 98562 273670
rect 99422 273670 99508 273730
rect 100672 273730 100732 274040
rect 101080 273730 101140 274040
rect 100672 273670 100770 273730
rect 98499 272916 98565 272917
rect 98499 272852 98500 272916
rect 98564 272852 98565 272916
rect 98499 272851 98565 272852
rect 99422 272237 99482 273670
rect 100710 272373 100770 273670
rect 101078 273670 101140 273730
rect 101760 273730 101820 274040
rect 102848 273730 102908 274040
rect 101760 273670 101874 273730
rect 100707 272372 100773 272373
rect 100707 272308 100708 272372
rect 100772 272308 100773 272372
rect 100707 272307 100773 272308
rect 99419 272236 99485 272237
rect 99419 272172 99420 272236
rect 99484 272172 99485 272236
rect 99419 272171 99485 272172
rect 98131 271828 98197 271829
rect 98131 271764 98132 271828
rect 98196 271764 98197 271828
rect 98131 271763 98197 271764
rect 95514 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 96134 260114
rect 95514 259794 96134 259878
rect 95514 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 96134 259794
rect 95514 252308 96134 259558
rect 99234 261954 99854 272000
rect 101078 271693 101138 273670
rect 101814 273189 101874 273670
rect 102734 273670 102908 273730
rect 103528 273730 103588 274040
rect 103936 273730 103996 274040
rect 103528 273670 103714 273730
rect 101811 273188 101877 273189
rect 101811 273124 101812 273188
rect 101876 273124 101877 273188
rect 101811 273123 101877 273124
rect 102734 271829 102794 273670
rect 102731 271828 102797 271829
rect 102731 271764 102732 271828
rect 102796 271764 102797 271828
rect 102731 271763 102797 271764
rect 101075 271692 101141 271693
rect 101075 271628 101076 271692
rect 101140 271628 101141 271692
rect 101075 271627 101141 271628
rect 99234 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 99854 261954
rect 99234 261634 99854 261718
rect 99234 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 99854 261634
rect 99234 252308 99854 261398
rect 102954 265674 103574 272000
rect 103654 271418 103714 273670
rect 103838 273670 103996 273730
rect 105296 273730 105356 274040
rect 105976 273730 106036 274040
rect 105296 273670 105370 273730
rect 103838 272781 103898 273670
rect 103835 272780 103901 272781
rect 103835 272716 103836 272780
rect 103900 272716 103901 272780
rect 103835 272715 103901 272716
rect 105310 271829 105370 273670
rect 105862 273670 106036 273730
rect 106384 273730 106444 274040
rect 107608 273866 107668 274040
rect 107518 273806 107668 273866
rect 106384 273670 106474 273730
rect 105307 271828 105373 271829
rect 105307 271764 105308 271828
rect 105372 271764 105373 271828
rect 105307 271763 105373 271764
rect 103835 271420 103901 271421
rect 103835 271418 103836 271420
rect 103654 271358 103836 271418
rect 103835 271356 103836 271358
rect 103900 271356 103901 271420
rect 103835 271355 103901 271356
rect 105862 271285 105922 273670
rect 105859 271284 105925 271285
rect 105859 271220 105860 271284
rect 105924 271220 105925 271284
rect 105859 271219 105925 271220
rect 106414 270877 106474 273670
rect 107518 271829 107578 273806
rect 108288 273730 108348 274040
rect 108696 273730 108756 274040
rect 109784 273730 109844 274040
rect 108254 273670 108348 273730
rect 108622 273670 108756 273730
rect 109542 273670 109844 273730
rect 111008 273730 111068 274040
rect 111144 273730 111204 274040
rect 112232 273730 112292 274040
rect 113320 273869 113380 274040
rect 113317 273868 113383 273869
rect 113317 273804 113318 273868
rect 113382 273804 113383 273868
rect 113317 273803 113383 273804
rect 113592 273730 113652 274040
rect 111008 273670 111074 273730
rect 111144 273670 111258 273730
rect 107515 271828 107581 271829
rect 107515 271764 107516 271828
rect 107580 271764 107581 271828
rect 107515 271763 107581 271764
rect 108254 271285 108314 273670
rect 108622 272509 108682 273670
rect 108619 272508 108685 272509
rect 108619 272444 108620 272508
rect 108684 272444 108685 272508
rect 108619 272443 108685 272444
rect 108251 271284 108317 271285
rect 108251 271220 108252 271284
rect 108316 271220 108317 271284
rect 108251 271219 108317 271220
rect 106411 270876 106477 270877
rect 106411 270812 106412 270876
rect 106476 270812 106477 270876
rect 106411 270811 106477 270812
rect 109542 270605 109602 273670
rect 109539 270604 109605 270605
rect 109539 270540 109540 270604
rect 109604 270540 109605 270604
rect 109539 270539 109605 270540
rect 102954 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 103574 265674
rect 102954 265354 103574 265438
rect 102954 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 103574 265354
rect 102954 252308 103574 265118
rect 109794 255454 110414 272000
rect 111014 271693 111074 273670
rect 111011 271692 111077 271693
rect 111011 271628 111012 271692
rect 111076 271628 111077 271692
rect 111011 271627 111077 271628
rect 111198 270605 111258 273670
rect 112118 273670 112292 273730
rect 113222 273670 113652 273730
rect 114408 273730 114468 274040
rect 115768 273730 115828 274040
rect 116040 273730 116100 274040
rect 116992 273730 117052 274040
rect 118080 273730 118140 274040
rect 118488 273730 118548 274040
rect 119168 273730 119228 274040
rect 120936 273730 120996 274040
rect 114408 273670 114570 273730
rect 115768 273670 115858 273730
rect 112118 271149 112178 273670
rect 113222 271421 113282 273670
rect 113219 271420 113285 271421
rect 113219 271356 113220 271420
rect 113284 271356 113285 271420
rect 113219 271355 113285 271356
rect 112115 271148 112181 271149
rect 112115 271084 112116 271148
rect 112180 271084 112181 271148
rect 112115 271083 112181 271084
rect 111195 270604 111261 270605
rect 111195 270540 111196 270604
rect 111260 270540 111261 270604
rect 111195 270539 111261 270540
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 252308 110414 254898
rect 113514 259174 114134 272000
rect 114510 271829 114570 273670
rect 114507 271828 114573 271829
rect 114507 271764 114508 271828
rect 114572 271764 114573 271828
rect 114507 271763 114573 271764
rect 115798 271013 115858 273670
rect 115982 273670 116100 273730
rect 116902 273670 117052 273730
rect 118006 273670 118140 273730
rect 118374 273670 118548 273730
rect 119110 273670 119228 273730
rect 120766 273670 120996 273730
rect 123520 273730 123580 274040
rect 125968 273730 126028 274040
rect 123520 273670 123586 273730
rect 115982 271557 116042 273670
rect 115979 271556 116045 271557
rect 115979 271492 115980 271556
rect 116044 271492 116045 271556
rect 115979 271491 116045 271492
rect 115795 271012 115861 271013
rect 115795 270948 115796 271012
rect 115860 270948 115861 271012
rect 115795 270947 115861 270948
rect 116902 270877 116962 273670
rect 118006 272645 118066 273670
rect 118003 272644 118069 272645
rect 118003 272580 118004 272644
rect 118068 272580 118069 272644
rect 118003 272579 118069 272580
rect 116899 270876 116965 270877
rect 116899 270812 116900 270876
rect 116964 270812 116965 270876
rect 116899 270811 116965 270812
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 252308 114134 258618
rect 117234 262894 117854 272000
rect 118374 271557 118434 273670
rect 118371 271556 118437 271557
rect 118371 271492 118372 271556
rect 118436 271492 118437 271556
rect 118371 271491 118437 271492
rect 119110 271285 119170 273670
rect 120766 271693 120826 273670
rect 120763 271692 120829 271693
rect 120763 271628 120764 271692
rect 120828 271628 120829 271692
rect 120763 271627 120829 271628
rect 119107 271284 119173 271285
rect 119107 271220 119108 271284
rect 119172 271220 119173 271284
rect 119107 271219 119173 271220
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 252308 117854 262338
rect 120954 266614 121574 272000
rect 123526 271829 123586 273670
rect 125918 273670 126028 273730
rect 128280 273730 128340 274040
rect 131000 273730 131060 274040
rect 133448 273733 133508 274040
rect 128280 273670 128738 273730
rect 125918 271829 125978 273670
rect 123523 271828 123589 271829
rect 123523 271764 123524 271828
rect 123588 271764 123589 271828
rect 123523 271763 123589 271764
rect 125915 271828 125981 271829
rect 125915 271764 125916 271828
rect 125980 271764 125981 271828
rect 125915 271763 125981 271764
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 252308 121574 266058
rect 127794 256394 128414 272000
rect 128678 271693 128738 273670
rect 130886 273670 131060 273730
rect 133445 273732 133511 273733
rect 130886 271829 130946 273670
rect 133445 273668 133446 273732
rect 133510 273668 133511 273732
rect 133445 273667 133511 273668
rect 135896 273597 135956 274040
rect 138480 273597 138540 274040
rect 140928 273597 140988 274040
rect 143512 273597 143572 274040
rect 145960 273597 146020 274040
rect 148544 273730 148604 274040
rect 150992 273730 151052 274040
rect 148544 273670 148610 273730
rect 135893 273596 135959 273597
rect 135893 273532 135894 273596
rect 135958 273532 135959 273596
rect 135893 273531 135959 273532
rect 138477 273596 138543 273597
rect 138477 273532 138478 273596
rect 138542 273532 138543 273596
rect 138477 273531 138543 273532
rect 140925 273596 140991 273597
rect 140925 273532 140926 273596
rect 140990 273532 140991 273596
rect 140925 273531 140991 273532
rect 143509 273596 143575 273597
rect 143509 273532 143510 273596
rect 143574 273532 143575 273596
rect 143509 273531 143575 273532
rect 145957 273596 146023 273597
rect 145957 273532 145958 273596
rect 146022 273532 146023 273596
rect 145957 273531 146023 273532
rect 130883 271828 130949 271829
rect 130883 271764 130884 271828
rect 130948 271764 130949 271828
rect 130883 271763 130949 271764
rect 128675 271692 128741 271693
rect 128675 271628 128676 271692
rect 128740 271628 128741 271692
rect 128675 271627 128741 271628
rect 127794 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 128414 256394
rect 127794 256074 128414 256158
rect 127794 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 128414 256074
rect 127794 252308 128414 255838
rect 131514 260114 132134 272000
rect 131514 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 132134 260114
rect 131514 259794 132134 259878
rect 131514 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 132134 259794
rect 131514 252308 132134 259558
rect 135234 261954 135854 272000
rect 135234 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 135854 261954
rect 135234 261634 135854 261718
rect 135234 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 135854 261634
rect 135234 252308 135854 261398
rect 138954 265674 139574 272000
rect 138954 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 139574 265674
rect 138954 265354 139574 265438
rect 138954 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 139574 265354
rect 138954 252308 139574 265118
rect 145794 255454 146414 272000
rect 148550 270877 148610 273670
rect 150942 273670 151052 273730
rect 153440 273730 153500 274040
rect 155888 273730 155948 274040
rect 158472 273730 158532 274040
rect 160920 273730 160980 274040
rect 153440 273670 154130 273730
rect 155888 273670 155970 273730
rect 158472 273670 158546 273730
rect 148547 270876 148613 270877
rect 148547 270812 148548 270876
rect 148612 270812 148613 270876
rect 148547 270811 148613 270812
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 252308 146414 254898
rect 149514 259174 150134 272000
rect 150942 271829 151002 273670
rect 150939 271828 151005 271829
rect 150939 271764 150940 271828
rect 151004 271764 151005 271828
rect 150939 271763 151005 271764
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 252308 150134 258618
rect 153234 262894 153854 272000
rect 154070 271829 154130 273670
rect 154067 271828 154133 271829
rect 154067 271764 154068 271828
rect 154132 271764 154133 271828
rect 154067 271763 154133 271764
rect 155910 271693 155970 273670
rect 155907 271692 155973 271693
rect 155907 271628 155908 271692
rect 155972 271628 155973 271692
rect 155907 271627 155973 271628
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 252308 153854 262338
rect 156954 266614 157574 272000
rect 158486 271829 158546 273670
rect 160878 273670 160980 273730
rect 163368 273730 163428 274040
rect 165952 273730 166012 274040
rect 183224 273730 183284 274040
rect 163368 273670 163514 273730
rect 165952 273670 166090 273730
rect 158483 271828 158549 271829
rect 158483 271764 158484 271828
rect 158548 271764 158549 271828
rect 158483 271763 158549 271764
rect 160878 271693 160938 273670
rect 163454 271693 163514 273670
rect 160875 271692 160941 271693
rect 160875 271628 160876 271692
rect 160940 271628 160941 271692
rect 160875 271627 160941 271628
rect 163451 271692 163517 271693
rect 163451 271628 163452 271692
rect 163516 271628 163517 271692
rect 163451 271627 163517 271628
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 252308 157574 266058
rect 163794 256394 164414 272000
rect 166030 271693 166090 273670
rect 183142 273670 183284 273730
rect 183360 273730 183420 274040
rect 183360 273670 183570 273730
rect 166027 271692 166093 271693
rect 166027 271628 166028 271692
rect 166092 271628 166093 271692
rect 166027 271627 166093 271628
rect 163794 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 164414 256394
rect 163794 256074 164414 256158
rect 163794 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 164414 256074
rect 163794 252308 164414 255838
rect 167514 260114 168134 272000
rect 167514 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 168134 260114
rect 167514 259794 168134 259878
rect 167514 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 168134 259794
rect 167514 252308 168134 259558
rect 171234 261954 171854 272000
rect 171234 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 171854 261954
rect 171234 261634 171854 261718
rect 171234 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 171854 261634
rect 171234 252308 171854 261398
rect 174954 265674 175574 272000
rect 174954 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 175574 265674
rect 174954 265354 175574 265438
rect 174954 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 175574 265354
rect 174954 252308 175574 265118
rect 181794 255454 182414 272000
rect 183142 271693 183202 273670
rect 183139 271692 183205 271693
rect 183139 271628 183140 271692
rect 183204 271628 183205 271692
rect 183139 271627 183205 271628
rect 183510 270605 183570 273670
rect 183507 270604 183573 270605
rect 183507 270540 183508 270604
rect 183572 270540 183573 270604
rect 183507 270539 183573 270540
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 179643 253332 179709 253333
rect 179643 253268 179644 253332
rect 179708 253268 179709 253332
rect 179643 253267 179709 253268
rect 178539 253196 178605 253197
rect 178539 253132 178540 253196
rect 178604 253132 178605 253196
rect 178539 253131 178605 253132
rect 178542 250610 178602 253131
rect 178464 250550 178602 250610
rect 179646 250610 179706 253267
rect 181794 252308 182414 254898
rect 185514 259174 186134 272000
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 252308 186134 258618
rect 189234 262894 189854 272000
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 252308 189854 262338
rect 192954 266614 193574 272000
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 190867 253196 190933 253197
rect 190867 253132 190868 253196
rect 190932 253132 190933 253196
rect 190867 253131 190933 253132
rect 190870 250610 190930 253131
rect 192954 252308 193574 266058
rect 179646 250550 179748 250610
rect 178464 250240 178524 250550
rect 179688 250240 179748 250550
rect 190840 250550 190930 250610
rect 190840 250240 190900 250550
rect 60272 237454 60620 237486
rect 60272 237218 60328 237454
rect 60564 237218 60620 237454
rect 60272 237134 60620 237218
rect 60272 236898 60328 237134
rect 60564 236898 60620 237134
rect 60272 236866 60620 236898
rect 196000 237454 196348 237486
rect 196000 237218 196056 237454
rect 196292 237218 196348 237454
rect 196000 237134 196348 237218
rect 196000 236898 196056 237134
rect 196292 236898 196348 237134
rect 196000 236866 196348 236898
rect 60952 219454 61300 219486
rect 60952 219218 61008 219454
rect 61244 219218 61300 219454
rect 60952 219134 61300 219218
rect 60952 218898 61008 219134
rect 61244 218898 61300 219134
rect 60952 218866 61300 218898
rect 195320 219454 195668 219486
rect 195320 219218 195376 219454
rect 195612 219218 195668 219454
rect 195320 219134 195668 219218
rect 195320 218898 195376 219134
rect 195612 218898 195668 219134
rect 195320 218866 195668 218898
rect 60272 201454 60620 201486
rect 60272 201218 60328 201454
rect 60564 201218 60620 201454
rect 60272 201134 60620 201218
rect 60272 200898 60328 201134
rect 60564 200898 60620 201134
rect 60272 200866 60620 200898
rect 196000 201454 196348 201486
rect 196000 201218 196056 201454
rect 196292 201218 196348 201454
rect 196000 201134 196348 201218
rect 196000 200898 196056 201134
rect 196292 200898 196348 201134
rect 196000 200866 196348 200898
rect 60952 183454 61300 183486
rect 60952 183218 61008 183454
rect 61244 183218 61300 183454
rect 60952 183134 61300 183218
rect 60952 182898 61008 183134
rect 61244 182898 61300 183134
rect 60952 182866 61300 182898
rect 195320 183454 195668 183486
rect 195320 183218 195376 183454
rect 195612 183218 195668 183454
rect 195320 183134 195668 183218
rect 195320 182898 195376 183134
rect 195612 182898 195668 183134
rect 195320 182866 195668 182898
rect 76056 166290 76116 167106
rect 76054 166230 76116 166290
rect 77144 166290 77204 167106
rect 78232 166290 78292 167106
rect 79592 166290 79652 167106
rect 80544 167010 80604 167106
rect 81768 167010 81828 167106
rect 83128 167010 83188 167106
rect 84216 167010 84276 167106
rect 85440 167010 85500 167106
rect 77144 166230 77218 166290
rect 78232 166230 78322 166290
rect 59514 152114 60134 165000
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 60134 152114
rect 59514 151794 60134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 60134 151794
rect 59514 145308 60134 151558
rect 63234 155834 63854 165000
rect 63234 155598 63266 155834
rect 63502 155598 63586 155834
rect 63822 155598 63854 155834
rect 63234 155514 63854 155598
rect 63234 155278 63266 155514
rect 63502 155278 63586 155514
rect 63822 155278 63854 155514
rect 63234 145308 63854 155278
rect 66954 157674 67574 165000
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 67574 157674
rect 66954 157354 67574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 67574 157354
rect 66954 145308 67574 157118
rect 73794 147454 74414 165000
rect 76054 164253 76114 166230
rect 77158 164389 77218 166230
rect 77155 164388 77221 164389
rect 77155 164324 77156 164388
rect 77220 164324 77221 164388
rect 77155 164323 77221 164324
rect 76051 164252 76117 164253
rect 76051 164188 76052 164252
rect 76116 164188 76117 164252
rect 76051 164187 76117 164188
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 145308 74414 146898
rect 77514 151174 78134 165000
rect 78262 164253 78322 166230
rect 79550 166230 79652 166290
rect 80470 166950 80604 167010
rect 81758 166950 81828 167010
rect 83046 166950 83188 167010
rect 84150 166950 84276 167010
rect 85438 166950 85500 167010
rect 86528 167010 86588 167106
rect 87616 167010 87676 167106
rect 88296 167010 88356 167106
rect 88704 167010 88764 167106
rect 90064 167010 90124 167106
rect 86528 166950 86602 167010
rect 87616 166950 87706 167010
rect 88296 166950 88442 167010
rect 88704 166950 88810 167010
rect 79550 164253 79610 166230
rect 80470 164253 80530 166950
rect 81758 165613 81818 166950
rect 81755 165612 81821 165613
rect 81755 165548 81756 165612
rect 81820 165548 81821 165612
rect 81755 165547 81821 165548
rect 78259 164252 78325 164253
rect 78259 164188 78260 164252
rect 78324 164188 78325 164252
rect 78259 164187 78325 164188
rect 79547 164252 79613 164253
rect 79547 164188 79548 164252
rect 79612 164188 79613 164252
rect 79547 164187 79613 164188
rect 80467 164252 80533 164253
rect 80467 164188 80468 164252
rect 80532 164188 80533 164252
rect 80467 164187 80533 164188
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 145308 78134 150618
rect 81234 154894 81854 165000
rect 83046 164253 83106 166950
rect 84150 164253 84210 166950
rect 85438 165613 85498 166950
rect 85435 165612 85501 165613
rect 85435 165548 85436 165612
rect 85500 165548 85501 165612
rect 85435 165547 85501 165548
rect 83043 164252 83109 164253
rect 83043 164188 83044 164252
rect 83108 164188 83109 164252
rect 83043 164187 83109 164188
rect 84147 164252 84213 164253
rect 84147 164188 84148 164252
rect 84212 164188 84213 164252
rect 84147 164187 84213 164188
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 145308 81854 154338
rect 84954 158614 85574 165000
rect 86542 164253 86602 166950
rect 87646 164253 87706 166950
rect 88382 164797 88442 166950
rect 88379 164796 88445 164797
rect 88379 164732 88380 164796
rect 88444 164732 88445 164796
rect 88379 164731 88445 164732
rect 88750 164253 88810 166950
rect 90038 166950 90124 167010
rect 90744 167010 90804 167106
rect 91288 167010 91348 167106
rect 92376 167010 92436 167106
rect 93464 167010 93524 167106
rect 90744 166950 90834 167010
rect 91288 166950 91386 167010
rect 92376 166950 92490 167010
rect 90038 164253 90098 166950
rect 90774 164797 90834 166950
rect 90771 164796 90837 164797
rect 90771 164732 90772 164796
rect 90836 164732 90837 164796
rect 90771 164731 90837 164732
rect 91326 164253 91386 166950
rect 92430 165613 92490 166950
rect 93350 166950 93524 167010
rect 93600 167010 93660 167106
rect 94552 167010 94612 167106
rect 95912 167010 95972 167106
rect 93600 166950 93778 167010
rect 92427 165612 92493 165613
rect 92427 165548 92428 165612
rect 92492 165548 92493 165612
rect 92427 165547 92493 165548
rect 86539 164252 86605 164253
rect 86539 164188 86540 164252
rect 86604 164188 86605 164252
rect 86539 164187 86605 164188
rect 87643 164252 87709 164253
rect 87643 164188 87644 164252
rect 87708 164188 87709 164252
rect 87643 164187 87709 164188
rect 88747 164252 88813 164253
rect 88747 164188 88748 164252
rect 88812 164188 88813 164252
rect 88747 164187 88813 164188
rect 90035 164252 90101 164253
rect 90035 164188 90036 164252
rect 90100 164188 90101 164252
rect 90035 164187 90101 164188
rect 91323 164252 91389 164253
rect 91323 164188 91324 164252
rect 91388 164188 91389 164252
rect 91323 164187 91389 164188
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 145308 85574 158058
rect 91794 148394 92414 165000
rect 93350 164253 93410 166950
rect 93718 166837 93778 166950
rect 94454 166950 94612 167010
rect 95742 166950 95972 167010
rect 96048 167010 96108 167106
rect 97000 167010 97060 167106
rect 98088 167010 98148 167106
rect 98496 167010 98556 167106
rect 99448 167010 99508 167106
rect 96048 166950 96170 167010
rect 97000 166950 97090 167010
rect 98088 166950 98194 167010
rect 98496 166950 98562 167010
rect 93715 166836 93781 166837
rect 93715 166772 93716 166836
rect 93780 166772 93781 166836
rect 93715 166771 93781 166772
rect 94454 164253 94514 166950
rect 95742 165613 95802 166950
rect 96110 166837 96170 166950
rect 96107 166836 96173 166837
rect 96107 166772 96108 166836
rect 96172 166772 96173 166836
rect 96107 166771 96173 166772
rect 95739 165612 95805 165613
rect 95739 165548 95740 165612
rect 95804 165548 95805 165612
rect 95739 165547 95805 165548
rect 93347 164252 93413 164253
rect 93347 164188 93348 164252
rect 93412 164188 93413 164252
rect 93347 164187 93413 164188
rect 94451 164252 94517 164253
rect 94451 164188 94452 164252
rect 94516 164188 94517 164252
rect 94451 164187 94517 164188
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 92414 148394
rect 91794 148074 92414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 92414 148074
rect 91794 145308 92414 147838
rect 95514 152114 96134 165000
rect 97030 164525 97090 166950
rect 97027 164524 97093 164525
rect 97027 164460 97028 164524
rect 97092 164460 97093 164524
rect 97027 164459 97093 164460
rect 98134 164253 98194 166950
rect 98502 166837 98562 166950
rect 99422 166950 99508 167010
rect 100672 167010 100732 167106
rect 101080 167010 101140 167106
rect 100672 166950 100770 167010
rect 98499 166836 98565 166837
rect 98499 166772 98500 166836
rect 98564 166772 98565 166836
rect 98499 166771 98565 166772
rect 99422 165613 99482 166950
rect 99419 165612 99485 165613
rect 99419 165548 99420 165612
rect 99484 165548 99485 165612
rect 99419 165547 99485 165548
rect 98131 164252 98197 164253
rect 98131 164188 98132 164252
rect 98196 164188 98197 164252
rect 98131 164187 98197 164188
rect 95514 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 96134 152114
rect 95514 151794 96134 151878
rect 95514 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 96134 151794
rect 95514 145308 96134 151558
rect 99234 155834 99854 165000
rect 100710 164253 100770 166950
rect 101078 166950 101140 167010
rect 101760 167010 101820 167106
rect 102848 167010 102908 167106
rect 103528 167010 103588 167106
rect 103936 167010 103996 167106
rect 101760 166950 101874 167010
rect 101078 166837 101138 166950
rect 101075 166836 101141 166837
rect 101075 166772 101076 166836
rect 101140 166772 101141 166836
rect 101075 166771 101141 166772
rect 101814 164389 101874 166950
rect 102734 166950 102908 167010
rect 103470 166950 103588 167010
rect 103838 166950 103996 167010
rect 105296 167010 105356 167106
rect 105976 167010 106036 167106
rect 105296 166950 105370 167010
rect 101811 164388 101877 164389
rect 101811 164324 101812 164388
rect 101876 164324 101877 164388
rect 101811 164323 101877 164324
rect 102734 164253 102794 166950
rect 103470 165613 103530 166950
rect 103467 165612 103533 165613
rect 103467 165548 103468 165612
rect 103532 165548 103533 165612
rect 103467 165547 103533 165548
rect 100707 164252 100773 164253
rect 100707 164188 100708 164252
rect 100772 164188 100773 164252
rect 100707 164187 100773 164188
rect 102731 164252 102797 164253
rect 102731 164188 102732 164252
rect 102796 164188 102797 164252
rect 102731 164187 102797 164188
rect 99234 155598 99266 155834
rect 99502 155598 99586 155834
rect 99822 155598 99854 155834
rect 99234 155514 99854 155598
rect 99234 155278 99266 155514
rect 99502 155278 99586 155514
rect 99822 155278 99854 155514
rect 99234 145308 99854 155278
rect 102954 157674 103574 165000
rect 103838 164389 103898 166950
rect 103835 164388 103901 164389
rect 103835 164324 103836 164388
rect 103900 164324 103901 164388
rect 103835 164323 103901 164324
rect 105310 164253 105370 166950
rect 105862 166950 106036 167010
rect 106384 167010 106444 167106
rect 107608 167010 107668 167106
rect 108288 167010 108348 167106
rect 108696 167010 108756 167106
rect 106384 166950 106474 167010
rect 105862 166837 105922 166950
rect 105859 166836 105925 166837
rect 105859 166772 105860 166836
rect 105924 166772 105925 166836
rect 105859 166771 105925 166772
rect 106414 164253 106474 166950
rect 107518 166950 107668 167010
rect 108254 166950 108348 167010
rect 108622 166950 108756 167010
rect 107518 164253 107578 166950
rect 108254 166837 108314 166950
rect 108251 166836 108317 166837
rect 108251 166772 108252 166836
rect 108316 166772 108317 166836
rect 108251 166771 108317 166772
rect 108622 164253 108682 166950
rect 109784 166290 109844 167106
rect 109726 166230 109844 166290
rect 111008 166290 111068 167106
rect 111144 166565 111204 167106
rect 111141 166564 111207 166565
rect 111141 166500 111142 166564
rect 111206 166500 111207 166564
rect 111141 166499 111207 166500
rect 112232 166290 112292 167106
rect 113320 166290 113380 167106
rect 113592 166290 113652 167106
rect 111008 166230 111074 166290
rect 109726 165613 109786 166230
rect 111014 165613 111074 166230
rect 112118 166230 112292 166290
rect 113222 166230 113380 166290
rect 113590 166230 113652 166290
rect 114408 166290 114468 167106
rect 115768 166290 115828 167106
rect 116040 166290 116100 167106
rect 116992 166565 117052 167106
rect 116989 166564 117055 166565
rect 116989 166500 116990 166564
rect 117054 166500 117055 166564
rect 116989 166499 117055 166500
rect 118080 166290 118140 167106
rect 118488 166290 118548 167106
rect 119168 166290 119228 167106
rect 114408 166230 114570 166290
rect 115768 166230 115858 166290
rect 109723 165612 109789 165613
rect 109723 165548 109724 165612
rect 109788 165548 109789 165612
rect 109723 165547 109789 165548
rect 111011 165612 111077 165613
rect 111011 165548 111012 165612
rect 111076 165548 111077 165612
rect 111011 165547 111077 165548
rect 105307 164252 105373 164253
rect 105307 164188 105308 164252
rect 105372 164188 105373 164252
rect 105307 164187 105373 164188
rect 106411 164252 106477 164253
rect 106411 164188 106412 164252
rect 106476 164188 106477 164252
rect 106411 164187 106477 164188
rect 107515 164252 107581 164253
rect 107515 164188 107516 164252
rect 107580 164188 107581 164252
rect 107515 164187 107581 164188
rect 108619 164252 108685 164253
rect 108619 164188 108620 164252
rect 108684 164188 108685 164252
rect 108619 164187 108685 164188
rect 102954 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 103574 157674
rect 102954 157354 103574 157438
rect 102954 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 103574 157354
rect 102954 145308 103574 157118
rect 109794 147454 110414 165000
rect 112118 164661 112178 166230
rect 112115 164660 112181 164661
rect 112115 164596 112116 164660
rect 112180 164596 112181 164660
rect 112115 164595 112181 164596
rect 113222 164525 113282 166230
rect 113590 165613 113650 166230
rect 113587 165612 113653 165613
rect 113587 165548 113588 165612
rect 113652 165548 113653 165612
rect 113587 165547 113653 165548
rect 113219 164524 113285 164525
rect 113219 164460 113220 164524
rect 113284 164460 113285 164524
rect 113219 164459 113285 164460
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 145308 110414 146898
rect 113514 151174 114134 165000
rect 114510 164933 114570 166230
rect 114507 164932 114573 164933
rect 114507 164868 114508 164932
rect 114572 164868 114573 164932
rect 114507 164867 114573 164868
rect 115798 164661 115858 166230
rect 115982 166230 116100 166290
rect 118006 166230 118140 166290
rect 118374 166230 118548 166290
rect 119110 166230 119228 166290
rect 120936 166290 120996 167106
rect 123520 166290 123580 167106
rect 125968 166290 126028 167106
rect 128280 167010 128340 167106
rect 131000 167010 131060 167106
rect 128280 166950 128554 167010
rect 128280 166910 128370 166950
rect 120936 166230 121010 166290
rect 123520 166230 123586 166290
rect 115982 165613 116042 166230
rect 118006 165613 118066 166230
rect 118374 165613 118434 166230
rect 115979 165612 116045 165613
rect 115979 165548 115980 165612
rect 116044 165548 116045 165612
rect 115979 165547 116045 165548
rect 118003 165612 118069 165613
rect 118003 165548 118004 165612
rect 118068 165548 118069 165612
rect 118003 165547 118069 165548
rect 118371 165612 118437 165613
rect 118371 165548 118372 165612
rect 118436 165548 118437 165612
rect 118371 165547 118437 165548
rect 119110 165069 119170 166230
rect 120950 165613 121010 166230
rect 123526 165613 123586 166230
rect 125918 166230 126028 166290
rect 125918 165613 125978 166230
rect 128494 165613 128554 166950
rect 130886 166950 131060 167010
rect 133448 167010 133508 167106
rect 135896 167010 135956 167106
rect 133448 166950 133522 167010
rect 130886 165613 130946 166950
rect 133462 165613 133522 166950
rect 135854 166950 135956 167010
rect 135854 165613 135914 166950
rect 138480 166837 138540 167106
rect 140928 166837 140988 167106
rect 143512 166837 143572 167106
rect 145960 166837 146020 167106
rect 148544 167010 148604 167106
rect 150992 167010 151052 167106
rect 153440 167010 153500 167106
rect 148544 166950 148610 167010
rect 138477 166836 138543 166837
rect 138477 166772 138478 166836
rect 138542 166772 138543 166836
rect 138477 166771 138543 166772
rect 140925 166836 140991 166837
rect 140925 166772 140926 166836
rect 140990 166772 140991 166836
rect 140925 166771 140991 166772
rect 143509 166836 143575 166837
rect 143509 166772 143510 166836
rect 143574 166772 143575 166836
rect 143509 166771 143575 166772
rect 145957 166836 146023 166837
rect 145957 166772 145958 166836
rect 146022 166772 146023 166836
rect 145957 166771 146023 166772
rect 148550 166565 148610 166950
rect 150942 166950 151052 167010
rect 153334 166950 153500 167010
rect 155888 167010 155948 167106
rect 155888 166950 155970 167010
rect 148547 166564 148613 166565
rect 148547 166500 148548 166564
rect 148612 166500 148613 166564
rect 148547 166499 148613 166500
rect 150942 165613 151002 166950
rect 153334 166429 153394 166950
rect 153331 166428 153397 166429
rect 153331 166364 153332 166428
rect 153396 166364 153397 166428
rect 153331 166363 153397 166364
rect 120947 165612 121013 165613
rect 120947 165548 120948 165612
rect 121012 165548 121013 165612
rect 120947 165547 121013 165548
rect 123523 165612 123589 165613
rect 123523 165548 123524 165612
rect 123588 165548 123589 165612
rect 123523 165547 123589 165548
rect 125915 165612 125981 165613
rect 125915 165548 125916 165612
rect 125980 165548 125981 165612
rect 125915 165547 125981 165548
rect 128491 165612 128557 165613
rect 128491 165548 128492 165612
rect 128556 165548 128557 165612
rect 128491 165547 128557 165548
rect 130883 165612 130949 165613
rect 130883 165548 130884 165612
rect 130948 165548 130949 165612
rect 130883 165547 130949 165548
rect 133459 165612 133525 165613
rect 133459 165548 133460 165612
rect 133524 165548 133525 165612
rect 133459 165547 133525 165548
rect 135851 165612 135917 165613
rect 135851 165548 135852 165612
rect 135916 165548 135917 165612
rect 135851 165547 135917 165548
rect 150939 165612 151005 165613
rect 150939 165548 150940 165612
rect 151004 165548 151005 165612
rect 150939 165547 151005 165548
rect 155910 165341 155970 166950
rect 158472 166290 158532 167106
rect 160920 166290 160980 167106
rect 163368 166701 163428 167106
rect 163365 166700 163431 166701
rect 163365 166636 163366 166700
rect 163430 166636 163431 166700
rect 163365 166635 163431 166636
rect 158472 166230 158546 166290
rect 158486 165477 158546 166230
rect 160878 166230 160980 166290
rect 165952 166290 166012 167106
rect 183224 167010 183284 167106
rect 183142 166950 183284 167010
rect 183360 167010 183420 167106
rect 183360 166950 183570 167010
rect 165952 166230 166090 166290
rect 158483 165476 158549 165477
rect 158483 165412 158484 165476
rect 158548 165412 158549 165476
rect 158483 165411 158549 165412
rect 155907 165340 155973 165341
rect 155907 165276 155908 165340
rect 155972 165276 155973 165340
rect 155907 165275 155973 165276
rect 160878 165205 160938 166230
rect 166030 165477 166090 166230
rect 183142 165613 183202 166950
rect 183510 165613 183570 166950
rect 196574 166429 196634 485419
rect 196758 273053 196818 485691
rect 197859 485348 197925 485349
rect 197859 485284 197860 485348
rect 197924 485284 197925 485348
rect 197859 485283 197925 485284
rect 196755 273052 196821 273053
rect 196755 272988 196756 273052
rect 196820 272988 196821 273052
rect 196755 272987 196821 272988
rect 196571 166428 196637 166429
rect 196571 166364 196572 166428
rect 196636 166364 196637 166428
rect 196571 166363 196637 166364
rect 183139 165612 183205 165613
rect 183139 165548 183140 165612
rect 183204 165548 183205 165612
rect 183139 165547 183205 165548
rect 183507 165612 183573 165613
rect 183507 165548 183508 165612
rect 183572 165548 183573 165612
rect 183507 165547 183573 165548
rect 166027 165476 166093 165477
rect 166027 165412 166028 165476
rect 166092 165412 166093 165476
rect 166027 165411 166093 165412
rect 160875 165204 160941 165205
rect 160875 165140 160876 165204
rect 160940 165140 160941 165204
rect 160875 165139 160941 165140
rect 119107 165068 119173 165069
rect 119107 165004 119108 165068
rect 119172 165004 119173 165068
rect 119107 165003 119173 165004
rect 115795 164660 115861 164661
rect 115795 164596 115796 164660
rect 115860 164596 115861 164660
rect 115795 164595 115861 164596
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 145308 114134 150618
rect 117234 154894 117854 165000
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 145308 117854 154338
rect 120954 158614 121574 165000
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 145308 121574 158058
rect 127794 148394 128414 165000
rect 127794 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 128414 148394
rect 127794 148074 128414 148158
rect 127794 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 128414 148074
rect 127794 145308 128414 147838
rect 131514 152114 132134 165000
rect 131514 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 132134 152114
rect 131514 151794 132134 151878
rect 131514 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 132134 151794
rect 131514 145308 132134 151558
rect 135234 155834 135854 165000
rect 135234 155598 135266 155834
rect 135502 155598 135586 155834
rect 135822 155598 135854 155834
rect 135234 155514 135854 155598
rect 135234 155278 135266 155514
rect 135502 155278 135586 155514
rect 135822 155278 135854 155514
rect 135234 145308 135854 155278
rect 138954 157674 139574 165000
rect 138954 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 139574 157674
rect 138954 157354 139574 157438
rect 138954 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 139574 157354
rect 138954 145308 139574 157118
rect 145794 147454 146414 165000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 145308 146414 146898
rect 149514 151174 150134 165000
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 145308 150134 150618
rect 153234 154894 153854 165000
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 145308 153854 154338
rect 156954 158614 157574 165000
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 145308 157574 158058
rect 163794 148394 164414 165000
rect 163794 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 164414 148394
rect 163794 148074 164414 148158
rect 163794 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 164414 148074
rect 163794 145308 164414 147838
rect 167514 152114 168134 165000
rect 167514 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 168134 152114
rect 167514 151794 168134 151878
rect 167514 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 168134 151794
rect 167514 145308 168134 151558
rect 171234 155834 171854 165000
rect 171234 155598 171266 155834
rect 171502 155598 171586 155834
rect 171822 155598 171854 155834
rect 171234 155514 171854 155598
rect 171234 155278 171266 155514
rect 171502 155278 171586 155514
rect 171822 155278 171854 155514
rect 171234 145308 171854 155278
rect 174954 157674 175574 165000
rect 174954 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 175574 157674
rect 174954 157354 175574 157438
rect 174954 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 175574 157354
rect 174954 145308 175574 157118
rect 181794 147454 182414 165000
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 145308 182414 146898
rect 185514 151174 186134 165000
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 145308 186134 150618
rect 189234 154894 189854 165000
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 145308 189854 154338
rect 192954 158614 193574 165000
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 145308 193574 158058
rect 178539 144940 178605 144941
rect 178539 144876 178540 144940
rect 178604 144876 178605 144940
rect 178539 144875 178605 144876
rect 179643 144940 179709 144941
rect 179643 144876 179644 144940
rect 179708 144876 179709 144940
rect 179643 144875 179709 144876
rect 190867 144940 190933 144941
rect 190867 144876 190868 144940
rect 190932 144876 190933 144940
rect 190867 144875 190933 144876
rect 178542 143850 178602 144875
rect 178464 143790 178602 143850
rect 179646 143850 179706 144875
rect 190870 143850 190930 144875
rect 179646 143790 179748 143850
rect 178464 143202 178524 143790
rect 179688 143202 179748 143790
rect 190840 143790 190930 143850
rect 190840 143202 190900 143790
rect 60272 129454 60620 129486
rect 60272 129218 60328 129454
rect 60564 129218 60620 129454
rect 60272 129134 60620 129218
rect 60272 128898 60328 129134
rect 60564 128898 60620 129134
rect 60272 128866 60620 128898
rect 196000 129454 196348 129486
rect 196000 129218 196056 129454
rect 196292 129218 196348 129454
rect 196000 129134 196348 129218
rect 196000 128898 196056 129134
rect 196292 128898 196348 129134
rect 196000 128866 196348 128898
rect 60952 111454 61300 111486
rect 60952 111218 61008 111454
rect 61244 111218 61300 111454
rect 60952 111134 61300 111218
rect 60952 110898 61008 111134
rect 61244 110898 61300 111134
rect 60952 110866 61300 110898
rect 195320 111454 195668 111486
rect 195320 111218 195376 111454
rect 195612 111218 195668 111454
rect 195320 111134 195668 111218
rect 195320 110898 195376 111134
rect 195612 110898 195668 111134
rect 195320 110866 195668 110898
rect 60272 93454 60620 93486
rect 60272 93218 60328 93454
rect 60564 93218 60620 93454
rect 60272 93134 60620 93218
rect 60272 92898 60328 93134
rect 60564 92898 60620 93134
rect 60272 92866 60620 92898
rect 196000 93454 196348 93486
rect 196000 93218 196056 93454
rect 196292 93218 196348 93454
rect 196000 93134 196348 93218
rect 196000 92898 196056 93134
rect 196292 92898 196348 93134
rect 196000 92866 196348 92898
rect 60952 75454 61300 75486
rect 60952 75218 61008 75454
rect 61244 75218 61300 75454
rect 60952 75134 61300 75218
rect 60952 74898 61008 75134
rect 61244 74898 61300 75134
rect 60952 74866 61300 74898
rect 195320 75454 195668 75486
rect 195320 75218 195376 75454
rect 195612 75218 195668 75454
rect 195320 75134 195668 75218
rect 195320 74898 195376 75134
rect 195612 74898 195668 75134
rect 195320 74866 195668 74898
rect 76056 59530 76116 60106
rect 77144 59805 77204 60106
rect 77141 59804 77207 59805
rect 77141 59740 77142 59804
rect 77206 59740 77207 59804
rect 77141 59739 77207 59740
rect 76054 59470 76116 59530
rect 78232 59530 78292 60106
rect 79592 59530 79652 60106
rect 80544 59530 80604 60106
rect 78232 59470 78322 59530
rect 59307 58716 59373 58717
rect 59307 58652 59308 58716
rect 59372 58652 59373 58716
rect 59307 58651 59373 58652
rect 59123 58444 59189 58445
rect 59123 58380 59124 58444
rect 59188 58380 59189 58444
rect 59123 58379 59189 58380
rect 58939 57084 59005 57085
rect 58939 57020 58940 57084
rect 59004 57020 59005 57084
rect 58939 57019 59005 57020
rect 57467 54772 57533 54773
rect 57467 54708 57468 54772
rect 57532 54708 57533 54772
rect 57467 54707 57533 54708
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 76054 57901 76114 59470
rect 76051 57900 76117 57901
rect 76051 57836 76052 57900
rect 76116 57836 76117 57900
rect 76051 57835 76117 57836
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 78262 57901 78322 59470
rect 79550 59470 79652 59530
rect 80470 59470 80604 59530
rect 81768 59530 81828 60106
rect 83128 59805 83188 60106
rect 83125 59804 83191 59805
rect 83125 59740 83126 59804
rect 83190 59740 83191 59804
rect 83125 59739 83191 59740
rect 84216 59530 84276 60106
rect 85440 59530 85500 60106
rect 81768 59470 82002 59530
rect 79550 57901 79610 59470
rect 80470 57901 80530 59470
rect 78259 57900 78325 57901
rect 78259 57836 78260 57900
rect 78324 57836 78325 57900
rect 78259 57835 78325 57836
rect 79547 57900 79613 57901
rect 79547 57836 79548 57900
rect 79612 57836 79613 57900
rect 79547 57835 79613 57836
rect 80467 57900 80533 57901
rect 80467 57836 80468 57900
rect 80532 57836 80533 57900
rect 80467 57835 80533 57836
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81942 57901 82002 59470
rect 83966 59470 84276 59530
rect 85438 59470 85500 59530
rect 86528 59530 86588 60106
rect 87616 59530 87676 60106
rect 88296 59530 88356 60106
rect 88704 59530 88764 60106
rect 90064 59530 90124 60106
rect 86528 59470 86602 59530
rect 87616 59470 87706 59530
rect 88296 59470 88442 59530
rect 88704 59470 88810 59530
rect 83966 58037 84026 59470
rect 85438 58173 85498 59470
rect 85435 58172 85501 58173
rect 85435 58108 85436 58172
rect 85500 58108 85501 58172
rect 85435 58107 85501 58108
rect 83963 58036 84029 58037
rect 83963 57972 83964 58036
rect 84028 57972 84029 58036
rect 83963 57971 84029 57972
rect 81939 57900 82005 57901
rect 81939 57836 81940 57900
rect 82004 57836 82005 57900
rect 81939 57835 82005 57836
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 86542 57901 86602 59470
rect 87646 57901 87706 59470
rect 86539 57900 86605 57901
rect 86539 57836 86540 57900
rect 86604 57836 86605 57900
rect 86539 57835 86605 57836
rect 87643 57900 87709 57901
rect 87643 57836 87644 57900
rect 87708 57836 87709 57900
rect 87643 57835 87709 57836
rect 88382 57221 88442 59470
rect 88750 57901 88810 59470
rect 90038 59470 90124 59530
rect 90744 59530 90804 60106
rect 91288 59530 91348 60106
rect 92376 59530 92436 60106
rect 93464 59530 93524 60106
rect 90744 59470 90834 59530
rect 91288 59470 91386 59530
rect 90038 57901 90098 59470
rect 90774 57901 90834 59470
rect 91326 57901 91386 59470
rect 92246 59470 92436 59530
rect 93350 59470 93524 59530
rect 93600 59530 93660 60106
rect 94552 59669 94612 60106
rect 94549 59668 94615 59669
rect 94549 59604 94550 59668
rect 94614 59604 94615 59668
rect 94549 59603 94615 59604
rect 95912 59533 95972 60106
rect 96048 59666 96108 60106
rect 97000 59669 97060 60106
rect 98088 59669 98148 60106
rect 96997 59668 97063 59669
rect 96048 59606 96354 59666
rect 95912 59532 95989 59533
rect 93600 59470 93778 59530
rect 95912 59470 95924 59532
rect 92246 58173 92306 59470
rect 92243 58172 92309 58173
rect 92243 58108 92244 58172
rect 92308 58108 92309 58172
rect 92243 58107 92309 58108
rect 88747 57900 88813 57901
rect 88747 57836 88748 57900
rect 88812 57836 88813 57900
rect 88747 57835 88813 57836
rect 90035 57900 90101 57901
rect 90035 57836 90036 57900
rect 90100 57836 90101 57900
rect 90035 57835 90101 57836
rect 90771 57900 90837 57901
rect 90771 57836 90772 57900
rect 90836 57836 90837 57900
rect 90771 57835 90837 57836
rect 91323 57900 91389 57901
rect 91323 57836 91324 57900
rect 91388 57836 91389 57900
rect 91323 57835 91389 57836
rect 91794 57454 92414 58000
rect 93350 57901 93410 59470
rect 93718 57901 93778 59470
rect 95923 59468 95924 59470
rect 95988 59468 95989 59532
rect 95923 59467 95989 59468
rect 93347 57900 93413 57901
rect 93347 57836 93348 57900
rect 93412 57836 93413 57900
rect 93347 57835 93413 57836
rect 93715 57900 93781 57901
rect 93715 57836 93716 57900
rect 93780 57836 93781 57900
rect 93715 57835 93781 57836
rect 88379 57220 88445 57221
rect 88379 57156 88380 57220
rect 88444 57156 88445 57220
rect 88379 57155 88445 57156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 96294 57085 96354 59606
rect 96997 59604 96998 59668
rect 97062 59604 97063 59668
rect 96997 59603 97063 59604
rect 98085 59668 98151 59669
rect 98085 59604 98086 59668
rect 98150 59604 98151 59668
rect 98085 59603 98151 59604
rect 98496 59530 98556 60106
rect 99448 59530 99508 60106
rect 100672 59669 100732 60106
rect 100672 59668 100773 59669
rect 100672 59606 100708 59668
rect 100707 59604 100708 59606
rect 100772 59604 100773 59668
rect 100707 59603 100773 59604
rect 101080 59530 101140 60106
rect 101760 59805 101820 60106
rect 101757 59804 101823 59805
rect 101757 59740 101758 59804
rect 101822 59740 101823 59804
rect 101757 59739 101823 59740
rect 102848 59669 102908 60106
rect 102845 59668 102911 59669
rect 102845 59604 102846 59668
rect 102910 59604 102911 59668
rect 102845 59603 102911 59604
rect 98496 59470 98562 59530
rect 98502 57357 98562 59470
rect 99422 59470 99508 59530
rect 101078 59470 101140 59530
rect 103528 59530 103588 60106
rect 103936 59805 103996 60106
rect 103933 59804 103999 59805
rect 103933 59740 103934 59804
rect 103998 59740 103999 59804
rect 103933 59739 103999 59740
rect 105296 59530 105356 60106
rect 105976 59669 106036 60106
rect 105973 59668 106039 59669
rect 105973 59604 105974 59668
rect 106038 59604 106039 59668
rect 105973 59603 106039 59604
rect 106384 59530 106444 60106
rect 107608 59805 107668 60106
rect 107605 59804 107671 59805
rect 107605 59740 107606 59804
rect 107670 59740 107671 59804
rect 107605 59739 107671 59740
rect 108288 59530 108348 60106
rect 108696 59669 108756 60106
rect 108693 59668 108759 59669
rect 108693 59604 108694 59668
rect 108758 59604 108759 59668
rect 108693 59603 108759 59604
rect 109784 59530 109844 60106
rect 103528 59470 103898 59530
rect 105296 59470 105370 59530
rect 106384 59470 106474 59530
rect 99422 58173 99482 59470
rect 101078 58445 101138 59470
rect 101075 58444 101141 58445
rect 101075 58380 101076 58444
rect 101140 58380 101141 58444
rect 101075 58379 101141 58380
rect 99419 58172 99485 58173
rect 99419 58108 99420 58172
rect 99484 58108 99485 58172
rect 99419 58107 99485 58108
rect 98499 57356 98565 57357
rect 98499 57292 98500 57356
rect 98564 57292 98565 57356
rect 98499 57291 98565 57292
rect 96291 57084 96357 57085
rect 96291 57020 96292 57084
rect 96356 57020 96357 57084
rect 96291 57019 96357 57020
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 103838 57221 103898 59470
rect 105310 57493 105370 59470
rect 106414 57629 106474 59470
rect 108254 59470 108348 59530
rect 109542 59470 109844 59530
rect 111008 59530 111068 60106
rect 111144 59530 111204 60106
rect 112232 59530 112292 60106
rect 113320 59530 113380 60106
rect 113592 59805 113652 60106
rect 113589 59804 113655 59805
rect 113589 59740 113590 59804
rect 113654 59740 113655 59804
rect 113589 59739 113655 59740
rect 114408 59530 114468 60106
rect 111008 59470 111074 59530
rect 111144 59470 111258 59530
rect 108254 58581 108314 59470
rect 108251 58580 108317 58581
rect 108251 58516 108252 58580
rect 108316 58516 108317 58580
rect 108251 58515 108317 58516
rect 109542 57901 109602 59470
rect 111014 59397 111074 59470
rect 111011 59396 111077 59397
rect 111011 59332 111012 59396
rect 111076 59332 111077 59396
rect 111011 59331 111077 59332
rect 109539 57900 109605 57901
rect 109539 57836 109540 57900
rect 109604 57836 109605 57900
rect 109539 57835 109605 57836
rect 106411 57628 106477 57629
rect 106411 57564 106412 57628
rect 106476 57564 106477 57628
rect 106411 57563 106477 57564
rect 105307 57492 105373 57493
rect 105307 57428 105308 57492
rect 105372 57428 105373 57492
rect 105307 57427 105373 57428
rect 103835 57220 103901 57221
rect 103835 57156 103836 57220
rect 103900 57156 103901 57220
rect 103835 57155 103901 57156
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 111198 57629 111258 59470
rect 112118 59470 112292 59530
rect 113222 59470 113380 59530
rect 114326 59470 114468 59530
rect 115768 59530 115828 60106
rect 116040 59530 116100 60106
rect 116992 59530 117052 60106
rect 118080 59530 118140 60106
rect 118488 59530 118548 60106
rect 119168 59530 119228 60106
rect 115768 59470 115858 59530
rect 112118 57901 112178 59470
rect 112115 57900 112181 57901
rect 112115 57836 112116 57900
rect 112180 57836 112181 57900
rect 112115 57835 112181 57836
rect 113222 57629 113282 59470
rect 111195 57628 111261 57629
rect 111195 57564 111196 57628
rect 111260 57564 111261 57628
rect 111195 57563 111261 57564
rect 113219 57628 113285 57629
rect 113219 57564 113220 57628
rect 113284 57564 113285 57628
rect 113219 57563 113285 57564
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 114326 57901 114386 59470
rect 114323 57900 114389 57901
rect 114323 57836 114324 57900
rect 114388 57836 114389 57900
rect 114323 57835 114389 57836
rect 115798 57629 115858 59470
rect 115982 59470 116100 59530
rect 116902 59470 117052 59530
rect 118006 59470 118140 59530
rect 118374 59470 118548 59530
rect 119110 59470 119228 59530
rect 120936 59530 120996 60106
rect 123520 59530 123580 60106
rect 125968 59530 126028 60106
rect 120936 59470 121010 59530
rect 123520 59470 123586 59530
rect 115982 57901 116042 59470
rect 116902 57901 116962 59470
rect 115979 57900 116045 57901
rect 115979 57836 115980 57900
rect 116044 57836 116045 57900
rect 115979 57835 116045 57836
rect 116899 57900 116965 57901
rect 116899 57836 116900 57900
rect 116964 57836 116965 57900
rect 116899 57835 116965 57836
rect 115795 57628 115861 57629
rect 115795 57564 115796 57628
rect 115860 57564 115861 57628
rect 115795 57563 115861 57564
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 118006 57765 118066 59470
rect 118003 57764 118069 57765
rect 118003 57700 118004 57764
rect 118068 57700 118069 57764
rect 118003 57699 118069 57700
rect 118374 56813 118434 59470
rect 119110 57629 119170 59470
rect 120950 58717 121010 59470
rect 120947 58716 121013 58717
rect 120947 58652 120948 58716
rect 121012 58652 121013 58716
rect 120947 58651 121013 58652
rect 119107 57628 119173 57629
rect 119107 57564 119108 57628
rect 119172 57564 119173 57628
rect 119107 57563 119173 57564
rect 118371 56812 118437 56813
rect 118371 56748 118372 56812
rect 118436 56748 118437 56812
rect 118371 56747 118437 56748
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 123526 57901 123586 59470
rect 125918 59470 126028 59530
rect 128280 59530 128340 60106
rect 131000 59530 131060 60106
rect 128280 59470 128370 59530
rect 125918 57901 125978 59470
rect 128310 58173 128370 59470
rect 130886 59470 131060 59530
rect 133448 59530 133508 60106
rect 135896 59530 135956 60106
rect 138480 59530 138540 60106
rect 140928 59530 140988 60106
rect 133448 59470 133522 59530
rect 128307 58172 128373 58173
rect 128307 58108 128308 58172
rect 128372 58108 128373 58172
rect 128307 58107 128373 58108
rect 123523 57900 123589 57901
rect 123523 57836 123524 57900
rect 123588 57836 123589 57900
rect 123523 57835 123589 57836
rect 125915 57900 125981 57901
rect 125915 57836 125916 57900
rect 125980 57836 125981 57900
rect 125915 57835 125981 57836
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 130886 57901 130946 59470
rect 130883 57900 130949 57901
rect 130883 57836 130884 57900
rect 130948 57836 130949 57900
rect 130883 57835 130949 57836
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 133462 57901 133522 59470
rect 135854 59470 135956 59530
rect 138430 59470 138540 59530
rect 140822 59470 140988 59530
rect 143512 59530 143572 60106
rect 145960 59530 146020 60106
rect 143512 59470 143642 59530
rect 135854 58853 135914 59470
rect 138430 58989 138490 59470
rect 140822 59125 140882 59470
rect 143582 59261 143642 59470
rect 145606 59470 146020 59530
rect 148544 59530 148604 60106
rect 150992 59530 151052 60106
rect 153440 59530 153500 60106
rect 148544 59470 148610 59530
rect 143579 59260 143645 59261
rect 143579 59196 143580 59260
rect 143644 59196 143645 59260
rect 143579 59195 143645 59196
rect 140819 59124 140885 59125
rect 140819 59060 140820 59124
rect 140884 59060 140885 59124
rect 140819 59059 140885 59060
rect 138427 58988 138493 58989
rect 138427 58924 138428 58988
rect 138492 58924 138493 58988
rect 138427 58923 138493 58924
rect 135851 58852 135917 58853
rect 135851 58788 135852 58852
rect 135916 58788 135917 58852
rect 135851 58787 135917 58788
rect 133459 57900 133525 57901
rect 133459 57836 133460 57900
rect 133524 57836 133525 57900
rect 133459 57835 133525 57836
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 145606 57901 145666 59470
rect 148550 59261 148610 59470
rect 150942 59470 151052 59530
rect 153334 59470 153500 59530
rect 155888 59530 155948 60106
rect 158472 59530 158532 60106
rect 160920 59530 160980 60106
rect 163368 59530 163428 60106
rect 165952 59530 166012 60106
rect 183224 59530 183284 60106
rect 155888 59470 155970 59530
rect 158472 59470 158546 59530
rect 150942 59261 151002 59470
rect 148547 59260 148613 59261
rect 148547 59196 148548 59260
rect 148612 59196 148613 59260
rect 148547 59195 148613 59196
rect 150939 59260 151005 59261
rect 150939 59196 150940 59260
rect 151004 59196 151005 59260
rect 150939 59195 151005 59196
rect 153334 58173 153394 59470
rect 153331 58172 153397 58173
rect 153331 58108 153332 58172
rect 153396 58108 153397 58172
rect 153331 58107 153397 58108
rect 145603 57900 145669 57901
rect 145603 57836 145604 57900
rect 145668 57836 145669 57900
rect 145603 57835 145669 57836
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 155910 57629 155970 59470
rect 155907 57628 155973 57629
rect 155907 57564 155908 57628
rect 155972 57564 155973 57628
rect 155907 57563 155973 57564
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 158486 56405 158546 59470
rect 160878 59470 160980 59530
rect 163270 59470 163428 59530
rect 165846 59470 166012 59530
rect 183142 59470 183284 59530
rect 183360 59530 183420 60106
rect 183360 59470 183570 59530
rect 160878 57629 160938 59470
rect 160875 57628 160941 57629
rect 160875 57564 160876 57628
rect 160940 57564 160941 57628
rect 160875 57563 160941 57564
rect 163270 56677 163330 59470
rect 163794 57454 164414 58000
rect 165846 57629 165906 59470
rect 165843 57628 165909 57629
rect 165843 57564 165844 57628
rect 165908 57564 165909 57628
rect 165843 57563 165909 57564
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163267 56676 163333 56677
rect 163267 56612 163268 56676
rect 163332 56612 163333 56676
rect 163267 56611 163333 56612
rect 158483 56404 158549 56405
rect 158483 56340 158484 56404
rect 158548 56340 158549 56404
rect 158483 56339 158549 56340
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 183142 57901 183202 59470
rect 183139 57900 183205 57901
rect 183139 57836 183140 57900
rect 183204 57836 183205 57900
rect 183139 57835 183205 57836
rect 183510 57765 183570 59470
rect 197862 58717 197922 485283
rect 198595 485212 198661 485213
rect 198595 485148 198596 485212
rect 198660 485148 198661 485212
rect 198595 485147 198661 485148
rect 198043 484940 198109 484941
rect 198043 484876 198044 484940
rect 198108 484876 198109 484940
rect 198043 484875 198109 484876
rect 198046 273189 198106 484875
rect 198411 484804 198477 484805
rect 198411 484740 198412 484804
rect 198476 484740 198477 484804
rect 198411 484739 198477 484740
rect 198043 273188 198109 273189
rect 198043 273124 198044 273188
rect 198108 273124 198109 273188
rect 198043 273123 198109 273124
rect 198414 59261 198474 484739
rect 198411 59260 198477 59261
rect 198411 59196 198412 59260
rect 198476 59196 198477 59260
rect 198411 59195 198477 59196
rect 198598 58853 198658 485147
rect 198963 478140 199029 478141
rect 198963 478076 198964 478140
rect 199028 478076 199029 478140
rect 198963 478075 199029 478076
rect 198779 466308 198845 466309
rect 198779 466244 198780 466308
rect 198844 466244 198845 466308
rect 198779 466243 198845 466244
rect 198782 165477 198842 466243
rect 198966 397490 199026 478075
rect 199794 472394 200414 486000
rect 202275 485620 202341 485621
rect 202275 485556 202276 485620
rect 202340 485556 202341 485620
rect 202275 485555 202341 485556
rect 200619 485076 200685 485077
rect 200619 485012 200620 485076
rect 200684 485012 200685 485076
rect 200619 485011 200685 485012
rect 199794 472158 199826 472394
rect 200062 472158 200146 472394
rect 200382 472158 200414 472394
rect 199794 472074 200414 472158
rect 199794 471838 199826 472074
rect 200062 471838 200146 472074
rect 200382 471838 200414 472074
rect 199515 469164 199581 469165
rect 199515 469100 199516 469164
rect 199580 469100 199581 469164
rect 199515 469099 199581 469100
rect 199147 464404 199213 464405
rect 199147 464340 199148 464404
rect 199212 464340 199213 464404
rect 199147 464339 199213 464340
rect 199150 398037 199210 464339
rect 199147 398036 199213 398037
rect 199147 397972 199148 398036
rect 199212 397972 199213 398036
rect 199147 397971 199213 397972
rect 198966 397430 199394 397490
rect 199147 396132 199213 396133
rect 199147 396068 199148 396132
rect 199212 396068 199213 396132
rect 199147 396067 199213 396068
rect 199150 377909 199210 396067
rect 199334 395861 199394 397430
rect 199331 395860 199397 395861
rect 199331 395796 199332 395860
rect 199396 395796 199397 395860
rect 199331 395795 199397 395796
rect 199147 377908 199213 377909
rect 199147 377844 199148 377908
rect 199212 377844 199213 377908
rect 199147 377843 199213 377844
rect 199334 371925 199394 395795
rect 199518 379405 199578 469099
rect 199794 453454 200414 471838
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199515 379404 199581 379405
rect 199515 379340 199516 379404
rect 199580 379340 199581 379404
rect 199515 379339 199581 379340
rect 199331 371924 199397 371925
rect 199331 371860 199332 371924
rect 199396 371860 199397 371924
rect 199331 371859 199397 371860
rect 199794 364394 200414 380898
rect 199794 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 200414 364394
rect 199794 364074 200414 364158
rect 199794 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 200414 364074
rect 199794 345454 200414 363838
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 256394 200414 272898
rect 199794 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 200414 256394
rect 199794 256074 200414 256158
rect 199794 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 200414 256074
rect 199794 237454 200414 255838
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 198779 165476 198845 165477
rect 198779 165412 198780 165476
rect 198844 165412 198845 165476
rect 198779 165411 198845 165412
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 148394 200414 164898
rect 199794 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 200414 148394
rect 199794 148074 200414 148158
rect 199794 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 200414 148074
rect 199794 129454 200414 147838
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 198595 58852 198661 58853
rect 198595 58788 198596 58852
rect 198660 58788 198661 58852
rect 198595 58787 198661 58788
rect 197859 58716 197925 58717
rect 197859 58652 197860 58716
rect 197924 58652 197925 58716
rect 197859 58651 197925 58652
rect 183507 57764 183573 57765
rect 183507 57700 183508 57764
rect 183572 57700 183573 57764
rect 183507 57699 183573 57700
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 92898
rect 200622 58581 200682 485011
rect 201355 484804 201421 484805
rect 201355 484740 201356 484804
rect 201420 484740 201421 484804
rect 201355 484739 201421 484740
rect 200803 484668 200869 484669
rect 200803 484604 200804 484668
rect 200868 484604 200869 484668
rect 200803 484603 200869 484604
rect 200806 59397 200866 484603
rect 200987 469028 201053 469029
rect 200987 468964 200988 469028
rect 201052 468964 201053 469028
rect 200987 468963 201053 468964
rect 200990 164797 201050 468963
rect 200987 164796 201053 164797
rect 200987 164732 200988 164796
rect 201052 164732 201053 164796
rect 200987 164731 201053 164732
rect 200803 59396 200869 59397
rect 200803 59332 200804 59396
rect 200868 59332 200869 59396
rect 200803 59331 200869 59332
rect 200619 58580 200685 58581
rect 200619 58516 200620 58580
rect 200684 58516 200685 58580
rect 200619 58515 200685 58516
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 201358 56269 201418 484739
rect 202091 472564 202157 472565
rect 202091 472500 202092 472564
rect 202156 472500 202157 472564
rect 202091 472499 202157 472500
rect 202094 57221 202154 472499
rect 202278 166973 202338 485555
rect 202643 484940 202709 484941
rect 202643 484876 202644 484940
rect 202708 484876 202709 484940
rect 202643 484875 202709 484876
rect 202459 471748 202525 471749
rect 202459 471684 202460 471748
rect 202524 471684 202525 471748
rect 202459 471683 202525 471684
rect 202275 166972 202341 166973
rect 202275 166908 202276 166972
rect 202340 166908 202341 166972
rect 202275 166907 202341 166908
rect 202462 166837 202522 471683
rect 202646 379541 202706 484875
rect 203195 476916 203261 476917
rect 203195 476852 203196 476916
rect 203260 476852 203261 476916
rect 203195 476851 203261 476852
rect 203011 468892 203077 468893
rect 203011 468828 203012 468892
rect 203076 468828 203077 468892
rect 203011 468827 203077 468828
rect 202643 379540 202709 379541
rect 202643 379476 202644 379540
rect 202708 379476 202709 379540
rect 202643 379475 202709 379476
rect 202459 166836 202525 166837
rect 202459 166772 202460 166836
rect 202524 166772 202525 166836
rect 202459 166771 202525 166772
rect 203014 166701 203074 468827
rect 203011 166700 203077 166701
rect 203011 166636 203012 166700
rect 203076 166636 203077 166700
rect 203011 166635 203077 166636
rect 203198 57493 203258 476851
rect 203514 476114 204134 486000
rect 205403 485212 205469 485213
rect 205403 485148 205404 485212
rect 205468 485148 205469 485212
rect 205403 485147 205469 485148
rect 204851 478140 204917 478141
rect 204851 478076 204852 478140
rect 204916 478076 204917 478140
rect 204851 478075 204917 478076
rect 203514 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 204134 476114
rect 203514 475794 204134 475878
rect 203514 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 204134 475794
rect 203514 457174 204134 475558
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 368114 204134 384618
rect 203514 367878 203546 368114
rect 203782 367878 203866 368114
rect 204102 367878 204134 368114
rect 203514 367794 204134 367878
rect 203514 367558 203546 367794
rect 203782 367558 203866 367794
rect 204102 367558 204134 367794
rect 203514 349174 204134 367558
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 260114 204134 276618
rect 203514 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 204134 260114
rect 203514 259794 204134 259878
rect 203514 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 204134 259794
rect 203514 241174 204134 259558
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 152114 204134 168618
rect 203514 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 204134 152114
rect 203514 151794 204134 151878
rect 203514 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 204134 151794
rect 203514 133174 204134 151558
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203195 57492 203261 57493
rect 203195 57428 203196 57492
rect 203260 57428 203261 57492
rect 203195 57427 203261 57428
rect 202091 57220 202157 57221
rect 202091 57156 202092 57220
rect 202156 57156 202157 57220
rect 202091 57155 202157 57156
rect 201355 56268 201421 56269
rect 201355 56204 201356 56268
rect 201420 56204 201421 56268
rect 201355 56203 201421 56204
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 204854 4045 204914 478075
rect 205219 472836 205285 472837
rect 205219 472772 205220 472836
rect 205284 472772 205285 472836
rect 205219 472771 205285 472772
rect 205035 469844 205101 469845
rect 205035 469780 205036 469844
rect 205100 469780 205101 469844
rect 205035 469779 205101 469780
rect 205038 57765 205098 469779
rect 205222 165477 205282 472771
rect 205406 411365 205466 485147
rect 205771 483852 205837 483853
rect 205771 483788 205772 483852
rect 205836 483788 205837 483852
rect 205771 483787 205837 483788
rect 205774 476130 205834 483787
rect 205590 476070 205834 476130
rect 205403 411364 205469 411365
rect 205403 411300 205404 411364
rect 205468 411300 205469 411364
rect 205403 411299 205469 411300
rect 205590 381037 205650 476070
rect 205587 381036 205653 381037
rect 205587 380972 205588 381036
rect 205652 380972 205653 381036
rect 205587 380971 205653 380972
rect 205219 165476 205285 165477
rect 205219 165412 205220 165476
rect 205284 165412 205285 165476
rect 205219 165411 205285 165412
rect 205035 57764 205101 57765
rect 205035 57700 205036 57764
rect 205100 57700 205101 57764
rect 205035 57699 205101 57700
rect 204851 4044 204917 4045
rect 204851 3980 204852 4044
rect 204916 3980 204917 4044
rect 204851 3979 204917 3980
rect 206142 3229 206202 486371
rect 206875 485212 206941 485213
rect 206875 485148 206876 485212
rect 206940 485148 206941 485212
rect 206875 485147 206941 485148
rect 206323 472700 206389 472701
rect 206323 472636 206324 472700
rect 206388 472636 206389 472700
rect 206323 472635 206389 472636
rect 206326 165341 206386 472635
rect 206323 165340 206389 165341
rect 206323 165276 206324 165340
rect 206388 165276 206389 165340
rect 206323 165275 206389 165276
rect 206878 59125 206938 485147
rect 207234 477954 207854 486000
rect 208899 485076 208965 485077
rect 208899 485012 208900 485076
rect 208964 485012 208965 485076
rect 208899 485011 208965 485012
rect 208347 479500 208413 479501
rect 208347 479436 208348 479500
rect 208412 479436 208413 479500
rect 208347 479435 208413 479436
rect 207234 477718 207266 477954
rect 207502 477718 207586 477954
rect 207822 477718 207854 477954
rect 207234 477634 207854 477718
rect 207234 477398 207266 477634
rect 207502 477398 207586 477634
rect 207822 477398 207854 477634
rect 207234 460894 207854 477398
rect 207979 471612 208045 471613
rect 207979 471548 207980 471612
rect 208044 471548 208045 471612
rect 207979 471547 208045 471548
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 369954 207854 388338
rect 207234 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 207854 369954
rect 207234 369634 207854 369718
rect 207234 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 207854 369634
rect 207234 352894 207854 369398
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 261954 207854 280338
rect 207234 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 207854 261954
rect 207234 261634 207854 261718
rect 207234 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 207854 261634
rect 207234 244894 207854 261398
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 155834 207854 172338
rect 207982 163981 208042 471547
rect 208163 468484 208229 468485
rect 208163 468420 208164 468484
rect 208228 468420 208229 468484
rect 208163 468419 208229 468420
rect 208166 165205 208226 468419
rect 208350 390693 208410 479435
rect 208347 390692 208413 390693
rect 208347 390628 208348 390692
rect 208412 390628 208413 390692
rect 208347 390627 208413 390628
rect 208902 375461 208962 485011
rect 209083 484804 209149 484805
rect 209083 484740 209084 484804
rect 209148 484740 209149 484804
rect 209083 484739 209149 484740
rect 209086 379541 209146 484739
rect 210954 481674 211574 486000
rect 212395 485756 212461 485757
rect 212395 485692 212396 485756
rect 212460 485692 212461 485756
rect 212395 485691 212461 485692
rect 211659 484668 211725 484669
rect 211659 484604 211660 484668
rect 211724 484604 211725 484668
rect 211659 484603 211725 484604
rect 210954 481438 210986 481674
rect 211222 481438 211306 481674
rect 211542 481438 211574 481674
rect 210954 481354 211574 481438
rect 210954 481118 210986 481354
rect 211222 481118 211306 481354
rect 211542 481118 211574 481354
rect 210371 479500 210437 479501
rect 210371 479436 210372 479500
rect 210436 479436 210437 479500
rect 210371 479435 210437 479436
rect 209819 478276 209885 478277
rect 209819 478212 209820 478276
rect 209884 478212 209885 478276
rect 209819 478211 209885 478212
rect 209083 379540 209149 379541
rect 209083 379476 209084 379540
rect 209148 379476 209149 379540
rect 209083 379475 209149 379476
rect 209822 375597 209882 478211
rect 210003 475556 210069 475557
rect 210003 475492 210004 475556
rect 210068 475492 210069 475556
rect 210003 475491 210069 475492
rect 209819 375596 209885 375597
rect 209819 375532 209820 375596
rect 209884 375532 209885 375596
rect 209819 375531 209885 375532
rect 210006 375461 210066 475491
rect 208899 375460 208965 375461
rect 208899 375396 208900 375460
rect 208964 375396 208965 375460
rect 208899 375395 208965 375396
rect 210003 375460 210069 375461
rect 210003 375396 210004 375460
rect 210068 375396 210069 375460
rect 210003 375395 210069 375396
rect 208163 165204 208229 165205
rect 208163 165140 208164 165204
rect 208228 165140 208229 165204
rect 208163 165139 208229 165140
rect 207979 163980 208045 163981
rect 207979 163916 207980 163980
rect 208044 163916 208045 163980
rect 207979 163915 208045 163916
rect 207234 155598 207266 155834
rect 207502 155598 207586 155834
rect 207822 155598 207854 155834
rect 207234 155514 207854 155598
rect 207234 155278 207266 155514
rect 207502 155278 207586 155514
rect 207822 155278 207854 155514
rect 207234 136894 207854 155278
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 206875 59124 206941 59125
rect 206875 59060 206876 59124
rect 206940 59060 206941 59124
rect 206875 59059 206941 59060
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 206139 3228 206205 3229
rect 206139 3164 206140 3228
rect 206204 3164 206205 3228
rect 206139 3163 206205 3164
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28338
rect 210374 3909 210434 479435
rect 210954 464614 211574 481118
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 373674 211574 392058
rect 211662 378181 211722 484603
rect 211659 378180 211725 378181
rect 211659 378116 211660 378180
rect 211724 378116 211725 378180
rect 211659 378115 211725 378116
rect 210954 373438 210986 373674
rect 211222 373438 211306 373674
rect 211542 373438 211574 373674
rect 210954 373354 211574 373438
rect 210954 373118 210986 373354
rect 211222 373118 211306 373354
rect 211542 373118 211574 373354
rect 210954 356614 211574 373118
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 265674 211574 284058
rect 210954 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 211574 265674
rect 210954 265354 211574 265438
rect 210954 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 211574 265354
rect 210954 248614 211574 265118
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 157674 211574 176058
rect 210954 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 211574 157674
rect 210954 157354 211574 157438
rect 210954 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 211574 157354
rect 210954 140614 211574 157118
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 212398 58989 212458 485691
rect 213683 485620 213749 485621
rect 213683 485556 213684 485620
rect 213748 485556 213749 485620
rect 213683 485555 213749 485556
rect 213131 483716 213197 483717
rect 213131 483652 213132 483716
rect 213196 483652 213197 483716
rect 213131 483651 213197 483652
rect 212395 58988 212461 58989
rect 212395 58924 212396 58988
rect 212460 58924 212461 58988
rect 212395 58923 212461 58924
rect 213134 57629 213194 483651
rect 213315 479636 213381 479637
rect 213315 479572 213316 479636
rect 213380 479572 213381 479636
rect 213315 479571 213381 479572
rect 213131 57628 213197 57629
rect 213131 57564 213132 57628
rect 213196 57564 213197 57628
rect 213131 57563 213197 57564
rect 213318 57357 213378 479571
rect 213499 468620 213565 468621
rect 213499 468556 213500 468620
rect 213564 468556 213565 468620
rect 213499 468555 213565 468556
rect 213502 166565 213562 468555
rect 213686 376821 213746 485555
rect 217547 485348 217613 485349
rect 217547 485284 217548 485348
rect 217612 485284 217613 485348
rect 217547 485283 217613 485284
rect 216995 484532 217061 484533
rect 216995 484468 216996 484532
rect 217060 484468 217061 484532
rect 216995 484467 217061 484468
rect 213867 482356 213933 482357
rect 213867 482292 213868 482356
rect 213932 482292 213933 482356
rect 213867 482291 213933 482292
rect 213683 376820 213749 376821
rect 213683 376756 213684 376820
rect 213748 376756 213749 376820
rect 213683 376755 213749 376756
rect 213870 375597 213930 482291
rect 215339 480996 215405 480997
rect 215339 480932 215340 480996
rect 215404 480932 215405 480996
rect 215339 480931 215405 480932
rect 214051 476780 214117 476781
rect 214051 476716 214052 476780
rect 214116 476716 214117 476780
rect 214051 476715 214117 476716
rect 213867 375596 213933 375597
rect 213867 375532 213868 375596
rect 213932 375532 213933 375596
rect 213867 375531 213933 375532
rect 214054 375461 214114 476715
rect 214419 474060 214485 474061
rect 214419 473996 214420 474060
rect 214484 473996 214485 474060
rect 214419 473995 214485 473996
rect 214051 375460 214117 375461
rect 214051 375396 214052 375460
rect 214116 375396 214117 375460
rect 214051 375395 214117 375396
rect 213499 166564 213565 166565
rect 213499 166500 213500 166564
rect 213564 166500 213565 166564
rect 213499 166499 213565 166500
rect 214422 68101 214482 473995
rect 214603 471204 214669 471205
rect 214603 471140 214604 471204
rect 214668 471140 214669 471204
rect 214603 471139 214669 471140
rect 214606 164117 214666 471139
rect 215342 273325 215402 480931
rect 215891 480860 215957 480861
rect 215891 480796 215892 480860
rect 215956 480796 215957 480860
rect 215891 480795 215957 480796
rect 215339 273324 215405 273325
rect 215339 273260 215340 273324
rect 215404 273260 215405 273324
rect 215339 273259 215405 273260
rect 214603 164116 214669 164117
rect 214603 164052 214604 164116
rect 214668 164052 214669 164116
rect 214603 164051 214669 164052
rect 214419 68100 214485 68101
rect 214419 68036 214420 68100
rect 214484 68036 214485 68100
rect 214419 68035 214485 68036
rect 213315 57356 213381 57357
rect 213315 57292 213316 57356
rect 213380 57292 213381 57356
rect 213315 57291 213381 57292
rect 215894 57085 215954 480795
rect 216075 475420 216141 475421
rect 216075 475356 216076 475420
rect 216140 475356 216141 475420
rect 216075 475355 216141 475356
rect 215891 57084 215957 57085
rect 215891 57020 215892 57084
rect 215956 57020 215957 57084
rect 215891 57019 215957 57020
rect 216078 56677 216138 475355
rect 216998 380493 217058 484467
rect 217179 479772 217245 479773
rect 217179 479708 217180 479772
rect 217244 479708 217245 479772
rect 217179 479707 217245 479708
rect 216627 380492 216693 380493
rect 216627 380428 216628 380492
rect 216692 380428 216693 380492
rect 216627 380427 216693 380428
rect 216995 380492 217061 380493
rect 216995 380428 216996 380492
rect 217060 380428 217061 380492
rect 216995 380427 217061 380428
rect 216630 377909 216690 380427
rect 216627 377908 216693 377909
rect 216627 377844 216628 377908
rect 216692 377844 216693 377908
rect 216627 377843 216693 377844
rect 217182 271557 217242 479707
rect 217363 471476 217429 471477
rect 217363 471412 217364 471476
rect 217428 471412 217429 471476
rect 217363 471411 217429 471412
rect 217366 273325 217426 471411
rect 217550 378045 217610 485283
rect 217794 471454 218414 486000
rect 219203 485212 219269 485213
rect 219203 485148 219204 485212
rect 219268 485148 219269 485212
rect 219203 485147 219269 485148
rect 219019 485076 219085 485077
rect 219019 485012 219020 485076
rect 219084 485012 219085 485076
rect 219019 485011 219085 485012
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 466308 218414 470898
rect 218651 467124 218717 467125
rect 218651 467060 218652 467124
rect 218716 467060 218717 467124
rect 218651 467059 218717 467060
rect 217547 378044 217613 378045
rect 217547 377980 217548 378044
rect 217612 377980 217613 378044
rect 217547 377979 217613 377980
rect 217547 374916 217613 374917
rect 217547 374852 217548 374916
rect 217612 374852 217613 374916
rect 217547 374851 217613 374852
rect 217363 273324 217429 273325
rect 217363 273260 217364 273324
rect 217428 273260 217429 273324
rect 217363 273259 217429 273260
rect 217179 271556 217245 271557
rect 217179 271492 217180 271556
rect 217244 271492 217245 271556
rect 217179 271491 217245 271492
rect 217550 269925 217610 374851
rect 217794 363454 218414 379000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 359308 218414 362898
rect 217547 269924 217613 269925
rect 217547 269860 217548 269924
rect 217612 269860 217613 269924
rect 217547 269859 217613 269860
rect 217179 268700 217245 268701
rect 217179 268636 217180 268700
rect 217244 268636 217245 268700
rect 217179 268635 217245 268636
rect 217182 162621 217242 268635
rect 217794 255454 218414 272000
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 252308 218414 254898
rect 218654 165613 218714 467059
rect 218651 165612 218717 165613
rect 218651 165548 218652 165612
rect 218716 165548 218717 165612
rect 218651 165547 218717 165548
rect 217179 162620 217245 162621
rect 217179 162556 217180 162620
rect 217244 162556 217245 162620
rect 217179 162555 217245 162556
rect 217182 161490 217242 162555
rect 217182 161430 217610 161490
rect 217363 148340 217429 148341
rect 217363 148276 217364 148340
rect 217428 148276 217429 148340
rect 217363 148275 217429 148276
rect 216075 56676 216141 56677
rect 216075 56612 216076 56676
rect 216140 56612 216141 56676
rect 216075 56611 216141 56612
rect 217366 56133 217426 148275
rect 217550 58445 217610 161430
rect 217794 147454 218414 165000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 145308 218414 146898
rect 219022 60621 219082 485011
rect 219019 60620 219085 60621
rect 219019 60556 219020 60620
rect 219084 60556 219085 60620
rect 219019 60555 219085 60556
rect 217547 58444 217613 58445
rect 217547 58380 217548 58444
rect 217612 58380 217613 58444
rect 217547 58379 217613 58380
rect 217363 56132 217429 56133
rect 217363 56068 217364 56132
rect 217428 56068 217429 56132
rect 217363 56067 217429 56068
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 210371 3908 210437 3909
rect 210371 3844 210372 3908
rect 210436 3844 210437 3908
rect 210371 3843 210437 3844
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 219206 56541 219266 485147
rect 219939 484532 220005 484533
rect 219939 484468 219940 484532
rect 220004 484468 220005 484532
rect 219939 484467 220005 484468
rect 219203 56540 219269 56541
rect 219203 56476 219204 56540
rect 219268 56476 219269 56540
rect 219203 56475 219269 56476
rect 219942 56405 220002 484467
rect 221514 475174 222134 486000
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 466308 222134 474618
rect 225234 478894 225854 486000
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 466308 225854 478338
rect 228954 482614 229574 486000
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 466308 229574 482058
rect 235794 472394 236414 486000
rect 235794 472158 235826 472394
rect 236062 472158 236146 472394
rect 236382 472158 236414 472394
rect 235794 472074 236414 472158
rect 235794 471838 235826 472074
rect 236062 471838 236146 472074
rect 236382 471838 236414 472074
rect 235794 466308 236414 471838
rect 239514 476114 240134 486000
rect 239514 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 240134 476114
rect 239514 475794 240134 475878
rect 239514 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 240134 475794
rect 239514 466308 240134 475558
rect 243234 477954 243854 486000
rect 243234 477718 243266 477954
rect 243502 477718 243586 477954
rect 243822 477718 243854 477954
rect 243234 477634 243854 477718
rect 243234 477398 243266 477634
rect 243502 477398 243586 477634
rect 243822 477398 243854 477634
rect 243234 466308 243854 477398
rect 246954 481674 247574 486000
rect 246954 481438 246986 481674
rect 247222 481438 247306 481674
rect 247542 481438 247574 481674
rect 246954 481354 247574 481438
rect 246954 481118 246986 481354
rect 247222 481118 247306 481354
rect 247542 481118 247574 481354
rect 246954 466308 247574 481118
rect 253794 471454 254414 486000
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 466308 254414 470898
rect 257514 475174 258134 486000
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 466308 258134 474618
rect 261234 478894 261854 486000
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 466308 261854 478338
rect 264954 482614 265574 486000
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 466308 265574 482058
rect 271794 472394 272414 486000
rect 271794 472158 271826 472394
rect 272062 472158 272146 472394
rect 272382 472158 272414 472394
rect 271794 472074 272414 472158
rect 271794 471838 271826 472074
rect 272062 471838 272146 472074
rect 272382 471838 272414 472074
rect 271794 466308 272414 471838
rect 275514 476114 276134 486000
rect 275514 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 275514 475794 276134 475878
rect 275514 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 275514 466308 276134 475558
rect 279234 477954 279854 486000
rect 279234 477718 279266 477954
rect 279502 477718 279586 477954
rect 279822 477718 279854 477954
rect 279234 477634 279854 477718
rect 279234 477398 279266 477634
rect 279502 477398 279586 477634
rect 279822 477398 279854 477634
rect 279234 466308 279854 477398
rect 282954 481674 283574 486000
rect 282954 481438 282986 481674
rect 283222 481438 283306 481674
rect 283542 481438 283574 481674
rect 282954 481354 283574 481438
rect 282954 481118 282986 481354
rect 283222 481118 283306 481354
rect 283542 481118 283574 481354
rect 282954 466308 283574 481118
rect 289794 471454 290414 486000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 466308 290414 470898
rect 293514 475174 294134 486000
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 466308 294134 474618
rect 297234 478894 297854 486000
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 466308 297854 478338
rect 300954 482614 301574 486000
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 466308 301574 482058
rect 307794 466308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 466308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 466308 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 635033 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 635033 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 635033 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 635033 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 635033 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 635033 348134 636618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 635033 351854 640338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 635033 355574 644058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 635033 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 635033 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 635033 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 635033 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 635033 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 635033 384134 636618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 635033 387854 640338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 635033 391574 644058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 635033 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 635033 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 635033 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 635033 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 635033 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 635033 420134 636618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 635033 423854 640338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 635033 427574 644058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 635033 434414 650898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 329208 615454 329528 615486
rect 329208 615218 329250 615454
rect 329486 615218 329528 615454
rect 329208 615134 329528 615218
rect 329208 614898 329250 615134
rect 329486 614898 329528 615134
rect 329208 614866 329528 614898
rect 359928 615454 360248 615486
rect 359928 615218 359970 615454
rect 360206 615218 360248 615454
rect 359928 615134 360248 615218
rect 359928 614898 359970 615134
rect 360206 614898 360248 615134
rect 359928 614866 360248 614898
rect 390648 615454 390968 615486
rect 390648 615218 390690 615454
rect 390926 615218 390968 615454
rect 390648 615134 390968 615218
rect 390648 614898 390690 615134
rect 390926 614898 390968 615134
rect 390648 614866 390968 614898
rect 421368 615454 421688 615486
rect 421368 615218 421410 615454
rect 421646 615218 421688 615454
rect 421368 615134 421688 615218
rect 421368 614898 421410 615134
rect 421646 614898 421688 615134
rect 421368 614866 421688 614898
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 344568 597454 344888 597486
rect 344568 597218 344610 597454
rect 344846 597218 344888 597454
rect 344568 597134 344888 597218
rect 344568 596898 344610 597134
rect 344846 596898 344888 597134
rect 344568 596866 344888 596898
rect 375288 597454 375608 597486
rect 375288 597218 375330 597454
rect 375566 597218 375608 597454
rect 375288 597134 375608 597218
rect 375288 596898 375330 597134
rect 375566 596898 375608 597134
rect 375288 596866 375608 596898
rect 406008 597454 406328 597486
rect 406008 597218 406050 597454
rect 406286 597218 406328 597454
rect 406008 597134 406328 597218
rect 406008 596898 406050 597134
rect 406286 596898 406328 597134
rect 406008 596866 406328 596898
rect 436139 594828 436205 594829
rect 436139 594764 436140 594828
rect 436204 594764 436205 594828
rect 436139 594763 436205 594764
rect 329208 579454 329528 579486
rect 329208 579218 329250 579454
rect 329486 579218 329528 579454
rect 329208 579134 329528 579218
rect 329208 578898 329250 579134
rect 329486 578898 329528 579134
rect 329208 578866 329528 578898
rect 359928 579454 360248 579486
rect 359928 579218 359970 579454
rect 360206 579218 360248 579454
rect 359928 579134 360248 579218
rect 359928 578898 359970 579134
rect 360206 578898 360248 579134
rect 359928 578866 360248 578898
rect 390648 579454 390968 579486
rect 390648 579218 390690 579454
rect 390926 579218 390968 579454
rect 390648 579134 390968 579218
rect 390648 578898 390690 579134
rect 390926 578898 390968 579134
rect 390648 578866 390968 578898
rect 421368 579454 421688 579486
rect 421368 579218 421410 579454
rect 421646 579218 421688 579454
rect 421368 579134 421688 579218
rect 421368 578898 421410 579134
rect 421646 578898 421688 579134
rect 421368 578866 421688 578898
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 344568 561454 344888 561486
rect 344568 561218 344610 561454
rect 344846 561218 344888 561454
rect 344568 561134 344888 561218
rect 344568 560898 344610 561134
rect 344846 560898 344888 561134
rect 344568 560866 344888 560898
rect 375288 561454 375608 561486
rect 375288 561218 375330 561454
rect 375566 561218 375608 561454
rect 375288 561134 375608 561218
rect 375288 560898 375330 561134
rect 375566 560898 375608 561134
rect 375288 560866 375608 560898
rect 406008 561454 406328 561486
rect 406008 561218 406050 561454
rect 406286 561218 406328 561454
rect 406008 561134 406328 561218
rect 406008 560898 406050 561134
rect 406286 560898 406328 561134
rect 406008 560866 406328 560898
rect 329208 543454 329528 543486
rect 329208 543218 329250 543454
rect 329486 543218 329528 543454
rect 329208 543134 329528 543218
rect 329208 542898 329250 543134
rect 329486 542898 329528 543134
rect 329208 542866 329528 542898
rect 359928 543454 360248 543486
rect 359928 543218 359970 543454
rect 360206 543218 360248 543454
rect 359928 543134 360248 543218
rect 359928 542898 359970 543134
rect 360206 542898 360248 543134
rect 359928 542866 360248 542898
rect 390648 543454 390968 543486
rect 390648 543218 390690 543454
rect 390926 543218 390968 543454
rect 390648 543134 390968 543218
rect 390648 542898 390690 543134
rect 390926 542898 390968 543134
rect 390648 542866 390968 542898
rect 421368 543454 421688 543486
rect 421368 543218 421410 543454
rect 421646 543218 421688 543454
rect 421368 543134 421688 543218
rect 421368 542898 421410 543134
rect 421646 542898 421688 543134
rect 421368 542866 421688 542898
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 344568 525454 344888 525486
rect 344568 525218 344610 525454
rect 344846 525218 344888 525454
rect 344568 525134 344888 525218
rect 344568 524898 344610 525134
rect 344846 524898 344888 525134
rect 344568 524866 344888 524898
rect 375288 525454 375608 525486
rect 375288 525218 375330 525454
rect 375566 525218 375608 525454
rect 375288 525134 375608 525218
rect 375288 524898 375330 525134
rect 375566 524898 375608 525134
rect 375288 524866 375608 524898
rect 406008 525454 406328 525486
rect 406008 525218 406050 525454
rect 406286 525218 406328 525454
rect 406008 525134 406328 525218
rect 406008 524898 406050 525134
rect 406286 524898 406328 525134
rect 406008 524866 406328 524898
rect 436142 522341 436202 594763
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 436139 522340 436205 522341
rect 436139 522276 436140 522340
rect 436204 522276 436205 522340
rect 436139 522275 436205 522276
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 466308 319574 500058
rect 325794 507454 326414 520000
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 466308 326414 470898
rect 329514 511174 330134 520000
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 466308 330134 474618
rect 333234 514894 333854 520000
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 466308 333854 478338
rect 336954 518614 337574 520000
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 466308 337574 482058
rect 343794 489454 344414 520000
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 338435 466580 338501 466581
rect 338435 466516 338436 466580
rect 338500 466516 338501 466580
rect 338435 466515 338501 466516
rect 339723 466580 339789 466581
rect 339723 466516 339724 466580
rect 339788 466516 339789 466580
rect 339723 466515 339789 466516
rect 338438 464810 338498 466515
rect 339726 464810 339786 466515
rect 343794 466308 344414 488898
rect 347514 493174 348134 520000
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 466308 348134 492618
rect 351234 496894 351854 520000
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350947 466580 351013 466581
rect 350947 466516 350948 466580
rect 351012 466516 351013 466580
rect 350947 466515 351013 466516
rect 350950 464810 351010 466515
rect 351234 466308 351854 496338
rect 354954 500614 355574 520000
rect 360883 516764 360949 516765
rect 360883 516700 360884 516764
rect 360948 516700 360949 516764
rect 360883 516699 360949 516700
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 466308 355574 500058
rect 357939 485756 358005 485757
rect 357939 485692 357940 485756
rect 358004 485692 358005 485756
rect 357939 485691 358005 485692
rect 356651 484940 356717 484941
rect 356651 484876 356652 484940
rect 356716 484876 356717 484940
rect 356651 484875 356717 484876
rect 338438 464750 338524 464810
rect 338464 464202 338524 464750
rect 339688 464750 339786 464810
rect 350840 464750 351010 464810
rect 339688 464202 339748 464750
rect 350840 464202 350900 464750
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 220952 399454 221300 399486
rect 220952 399218 221008 399454
rect 221244 399218 221300 399454
rect 220952 399134 221300 399218
rect 220952 398898 221008 399134
rect 221244 398898 221300 399134
rect 220952 398866 221300 398898
rect 355320 399454 355668 399486
rect 355320 399218 355376 399454
rect 355612 399218 355668 399454
rect 355320 399134 355668 399218
rect 355320 398898 355376 399134
rect 355612 398898 355668 399134
rect 355320 398866 355668 398898
rect 236056 380765 236116 381106
rect 237144 380765 237204 381106
rect 236053 380764 236119 380765
rect 236053 380700 236054 380764
rect 236118 380700 236119 380764
rect 236053 380699 236119 380700
rect 237141 380764 237207 380765
rect 237141 380700 237142 380764
rect 237206 380700 237207 380764
rect 237141 380699 237207 380700
rect 238232 380490 238292 381106
rect 239592 380490 239652 381106
rect 238158 380430 238292 380490
rect 239262 380430 239652 380490
rect 240544 380490 240604 381106
rect 241768 380490 241828 381106
rect 243128 380765 243188 381106
rect 243125 380764 243191 380765
rect 243125 380700 243126 380764
rect 243190 380700 243191 380764
rect 243125 380699 243191 380700
rect 244216 380490 244276 381106
rect 245440 380765 245500 381106
rect 245437 380764 245503 380765
rect 245437 380700 245438 380764
rect 245502 380700 245503 380764
rect 245437 380699 245503 380700
rect 246528 380490 246588 381106
rect 247616 380490 247676 381106
rect 248296 380490 248356 381106
rect 248704 380490 248764 381106
rect 240544 380430 240610 380490
rect 241768 380430 241898 380490
rect 244216 380430 244290 380490
rect 221514 367174 222134 379000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 359308 222134 366618
rect 225234 370894 225854 379000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 359308 225854 370338
rect 228954 374614 229574 379000
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 359308 229574 374058
rect 235794 364394 236414 379000
rect 238158 378725 238218 380430
rect 239262 379133 239322 380430
rect 239259 379132 239325 379133
rect 239259 379068 239260 379132
rect 239324 379068 239325 379132
rect 239259 379067 239325 379068
rect 238155 378724 238221 378725
rect 238155 378660 238156 378724
rect 238220 378660 238221 378724
rect 238155 378659 238221 378660
rect 235794 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 236414 364394
rect 235794 364074 236414 364158
rect 235794 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 236414 364074
rect 235794 359308 236414 363838
rect 239514 368114 240134 379000
rect 240550 378453 240610 380430
rect 241467 378996 241533 378997
rect 241467 378932 241468 378996
rect 241532 378932 241533 378996
rect 241467 378931 241533 378932
rect 241470 378453 241530 378931
rect 241838 378861 241898 380430
rect 241835 378860 241901 378861
rect 241835 378796 241836 378860
rect 241900 378796 241901 378860
rect 241835 378795 241901 378796
rect 241838 378453 241898 378795
rect 240547 378452 240613 378453
rect 240547 378388 240548 378452
rect 240612 378388 240613 378452
rect 240547 378387 240613 378388
rect 241467 378452 241533 378453
rect 241467 378388 241468 378452
rect 241532 378388 241533 378452
rect 241467 378387 241533 378388
rect 241835 378452 241901 378453
rect 241835 378388 241836 378452
rect 241900 378388 241901 378452
rect 241835 378387 241901 378388
rect 239514 367878 239546 368114
rect 239782 367878 239866 368114
rect 240102 367878 240134 368114
rect 239514 367794 240134 367878
rect 239514 367558 239546 367794
rect 239782 367558 239866 367794
rect 240102 367558 240134 367794
rect 239514 359308 240134 367558
rect 243234 369954 243854 379000
rect 244230 378317 244290 380430
rect 246438 380430 246588 380490
rect 247542 380430 247676 380490
rect 248278 380430 248356 380490
rect 248646 380430 248764 380490
rect 250064 380490 250124 381106
rect 250744 380490 250804 381106
rect 251288 380490 251348 381106
rect 252376 380490 252436 381106
rect 253464 380490 253524 381106
rect 250064 380430 250178 380490
rect 246438 379405 246498 380430
rect 247542 379405 247602 380430
rect 246435 379404 246501 379405
rect 246435 379340 246436 379404
rect 246500 379340 246501 379404
rect 246435 379339 246501 379340
rect 247539 379404 247605 379405
rect 247539 379340 247540 379404
rect 247604 379340 247605 379404
rect 247539 379339 247605 379340
rect 244227 378316 244293 378317
rect 244227 378252 244228 378316
rect 244292 378252 244293 378316
rect 244227 378251 244293 378252
rect 243234 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 243854 369954
rect 243234 369634 243854 369718
rect 243234 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 243854 369634
rect 243234 359308 243854 369398
rect 246954 373674 247574 379000
rect 248278 378861 248338 380430
rect 248646 379405 248706 380430
rect 250118 379405 250178 380430
rect 250670 380430 250804 380490
rect 251222 380430 251348 380490
rect 252326 380430 252436 380490
rect 253430 380430 253524 380490
rect 253600 380490 253660 381106
rect 254552 380629 254612 381106
rect 255912 380629 255972 381106
rect 256048 380765 256108 381106
rect 256045 380764 256111 380765
rect 256045 380700 256046 380764
rect 256110 380700 256111 380764
rect 256045 380699 256111 380700
rect 257000 380629 257060 381106
rect 254549 380628 254615 380629
rect 254549 380564 254550 380628
rect 254614 380564 254615 380628
rect 254549 380563 254615 380564
rect 255909 380628 255975 380629
rect 255909 380564 255910 380628
rect 255974 380564 255975 380628
rect 255909 380563 255975 380564
rect 256997 380628 257063 380629
rect 256997 380564 256998 380628
rect 257062 380564 257063 380628
rect 256997 380563 257063 380564
rect 258088 380490 258148 381106
rect 258496 380490 258556 381106
rect 259448 380629 259508 381106
rect 260672 380629 260732 381106
rect 259445 380628 259511 380629
rect 259445 380564 259446 380628
rect 259510 380564 259511 380628
rect 259445 380563 259511 380564
rect 260669 380628 260735 380629
rect 260669 380564 260670 380628
rect 260734 380564 260735 380628
rect 260669 380563 260735 380564
rect 261080 380490 261140 381106
rect 261760 380490 261820 381106
rect 262848 380490 262908 381106
rect 253600 380430 253674 380490
rect 248643 379404 248709 379405
rect 248643 379340 248644 379404
rect 248708 379340 248709 379404
rect 248643 379339 248709 379340
rect 250115 379404 250181 379405
rect 250115 379340 250116 379404
rect 250180 379340 250181 379404
rect 250115 379339 250181 379340
rect 248275 378860 248341 378861
rect 248275 378796 248276 378860
rect 248340 378796 248341 378860
rect 248275 378795 248341 378796
rect 250670 378317 250730 380430
rect 251222 379405 251282 380430
rect 252326 379405 252386 380430
rect 253430 379405 253490 380430
rect 251219 379404 251285 379405
rect 251219 379340 251220 379404
rect 251284 379340 251285 379404
rect 251219 379339 251285 379340
rect 252323 379404 252389 379405
rect 252323 379340 252324 379404
rect 252388 379340 252389 379404
rect 252323 379339 252389 379340
rect 253427 379404 253493 379405
rect 253427 379340 253428 379404
rect 253492 379340 253493 379404
rect 253427 379339 253493 379340
rect 253614 378589 253674 380430
rect 258030 380430 258148 380490
rect 258398 380430 258556 380490
rect 260974 380430 261140 380490
rect 261710 380430 261820 380490
rect 262814 380430 262908 380490
rect 263528 380490 263588 381106
rect 263936 380901 263996 381106
rect 263933 380900 263999 380901
rect 263933 380836 263934 380900
rect 263998 380836 263999 380900
rect 263933 380835 263999 380836
rect 265296 380629 265356 381106
rect 265293 380628 265359 380629
rect 265293 380564 265294 380628
rect 265358 380564 265359 380628
rect 265293 380563 265359 380564
rect 265976 380490 266036 381106
rect 266384 380490 266444 381106
rect 267608 380490 267668 381106
rect 263528 380430 263610 380490
rect 258030 379530 258090 380430
rect 257846 379470 258090 379530
rect 257846 379405 257906 379470
rect 257843 379404 257909 379405
rect 257843 379340 257844 379404
rect 257908 379340 257909 379404
rect 257843 379339 257909 379340
rect 253611 378588 253677 378589
rect 253611 378524 253612 378588
rect 253676 378524 253677 378588
rect 253611 378523 253677 378524
rect 250667 378316 250733 378317
rect 250667 378252 250668 378316
rect 250732 378252 250733 378316
rect 250667 378251 250733 378252
rect 246954 373438 246986 373674
rect 247222 373438 247306 373674
rect 247542 373438 247574 373674
rect 246954 373354 247574 373438
rect 246954 373118 246986 373354
rect 247222 373118 247306 373354
rect 247542 373118 247574 373354
rect 246954 359308 247574 373118
rect 253794 363454 254414 379000
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 359308 254414 362898
rect 257514 367174 258134 379000
rect 258398 378589 258458 380430
rect 260974 378589 261034 380430
rect 261710 379405 261770 380430
rect 261707 379404 261773 379405
rect 261707 379340 261708 379404
rect 261772 379340 261773 379404
rect 261707 379339 261773 379340
rect 258395 378588 258461 378589
rect 258395 378524 258396 378588
rect 258460 378524 258461 378588
rect 258395 378523 258461 378524
rect 260971 378588 261037 378589
rect 260971 378524 260972 378588
rect 261036 378524 261037 378588
rect 260971 378523 261037 378524
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 359308 258134 366618
rect 261234 370894 261854 379000
rect 262814 378317 262874 380430
rect 263550 378589 263610 380430
rect 265942 380430 266036 380490
rect 266310 380430 266444 380490
rect 267598 380430 267668 380490
rect 268288 380490 268348 381106
rect 268696 380490 268756 381106
rect 269784 380765 269844 381106
rect 269781 380764 269847 380765
rect 269781 380700 269782 380764
rect 269846 380700 269847 380764
rect 269781 380699 269847 380700
rect 271008 380629 271068 381106
rect 271005 380628 271071 380629
rect 271005 380564 271006 380628
rect 271070 380564 271071 380628
rect 271005 380563 271071 380564
rect 271144 380490 271204 381106
rect 272232 380490 272292 381106
rect 273320 380490 273380 381106
rect 273592 380490 273652 381106
rect 274408 380490 274468 381106
rect 275768 380490 275828 381106
rect 268288 380430 268394 380490
rect 268696 380430 268762 380490
rect 263547 378588 263613 378589
rect 263547 378524 263548 378588
rect 263612 378524 263613 378588
rect 263547 378523 263613 378524
rect 262811 378316 262877 378317
rect 262811 378252 262812 378316
rect 262876 378252 262877 378316
rect 262811 378251 262877 378252
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 359308 261854 370338
rect 264954 374614 265574 379000
rect 265942 378589 266002 380430
rect 265939 378588 266005 378589
rect 265939 378524 265940 378588
rect 266004 378524 266005 378588
rect 265939 378523 266005 378524
rect 266310 378317 266370 380430
rect 267598 378317 267658 380430
rect 268334 378589 268394 380430
rect 268702 379405 268762 380430
rect 271094 380430 271204 380490
rect 272198 380430 272292 380490
rect 273302 380430 273380 380490
rect 273486 380430 273652 380490
rect 274406 380430 274468 380490
rect 275694 380430 275828 380490
rect 276040 380490 276100 381106
rect 276992 380490 277052 381106
rect 276040 380430 276122 380490
rect 271094 379405 271154 380430
rect 272198 379405 272258 380430
rect 273302 379405 273362 380430
rect 268699 379404 268765 379405
rect 268699 379340 268700 379404
rect 268764 379340 268765 379404
rect 268699 379339 268765 379340
rect 271091 379404 271157 379405
rect 271091 379340 271092 379404
rect 271156 379340 271157 379404
rect 271091 379339 271157 379340
rect 272195 379404 272261 379405
rect 272195 379340 272196 379404
rect 272260 379340 272261 379404
rect 272195 379339 272261 379340
rect 273299 379404 273365 379405
rect 273299 379340 273300 379404
rect 273364 379340 273365 379404
rect 273299 379339 273365 379340
rect 268331 378588 268397 378589
rect 268331 378524 268332 378588
rect 268396 378524 268397 378588
rect 268331 378523 268397 378524
rect 266307 378316 266373 378317
rect 266307 378252 266308 378316
rect 266372 378252 266373 378316
rect 266307 378251 266373 378252
rect 267595 378316 267661 378317
rect 267595 378252 267596 378316
rect 267660 378252 267661 378316
rect 267595 378251 267661 378252
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 359308 265574 374058
rect 271794 364394 272414 379000
rect 273486 378589 273546 380430
rect 274406 379405 274466 380430
rect 275694 379405 275754 380430
rect 276062 379405 276122 380430
rect 276982 380430 277052 380490
rect 278080 380490 278140 381106
rect 278488 380490 278548 381106
rect 278080 380430 278146 380490
rect 276982 379405 277042 380430
rect 278086 379405 278146 380430
rect 278454 380430 278548 380490
rect 279168 380490 279228 381106
rect 280936 380490 280996 381106
rect 283520 380490 283580 381106
rect 279168 380430 279250 380490
rect 274403 379404 274469 379405
rect 274403 379340 274404 379404
rect 274468 379340 274469 379404
rect 274403 379339 274469 379340
rect 275691 379404 275757 379405
rect 275691 379340 275692 379404
rect 275756 379340 275757 379404
rect 275691 379339 275757 379340
rect 276059 379404 276125 379405
rect 276059 379340 276060 379404
rect 276124 379340 276125 379404
rect 276059 379339 276125 379340
rect 276979 379404 277045 379405
rect 276979 379340 276980 379404
rect 277044 379340 277045 379404
rect 276979 379339 277045 379340
rect 278083 379404 278149 379405
rect 278083 379340 278084 379404
rect 278148 379340 278149 379404
rect 278083 379339 278149 379340
rect 278454 379269 278514 380430
rect 279190 379269 279250 380430
rect 280846 380430 280996 380490
rect 283422 380430 283580 380490
rect 285968 380490 286028 381106
rect 288280 380490 288340 381106
rect 291000 380490 291060 381106
rect 293448 380490 293508 381106
rect 285968 380430 286058 380490
rect 280846 379269 280906 380430
rect 283422 379269 283482 380430
rect 285998 379405 286058 380430
rect 288206 380430 288340 380490
rect 290966 380430 291060 380490
rect 293358 380430 293508 380490
rect 295896 380490 295956 381106
rect 298480 380490 298540 381106
rect 300928 380490 300988 381106
rect 303512 380490 303572 381106
rect 305960 380490 306020 381106
rect 295896 380430 295994 380490
rect 298480 380430 298570 380490
rect 288206 379405 288266 380430
rect 290966 379405 291026 380430
rect 293358 379405 293418 380430
rect 295934 379405 295994 380430
rect 298510 379405 298570 380430
rect 300902 380430 300988 380490
rect 303478 380430 303572 380490
rect 305870 380430 306020 380490
rect 308544 380490 308604 381106
rect 310992 380490 311052 381106
rect 313440 380490 313500 381106
rect 315888 380490 315948 381106
rect 318472 380490 318532 381106
rect 308544 380430 308690 380490
rect 310992 380430 311082 380490
rect 300902 379405 300962 380430
rect 303478 379405 303538 380430
rect 305870 379405 305930 380430
rect 285995 379404 286061 379405
rect 285995 379340 285996 379404
rect 286060 379340 286061 379404
rect 285995 379339 286061 379340
rect 288203 379404 288269 379405
rect 288203 379340 288204 379404
rect 288268 379340 288269 379404
rect 288203 379339 288269 379340
rect 290963 379404 291029 379405
rect 290963 379340 290964 379404
rect 291028 379340 291029 379404
rect 290963 379339 291029 379340
rect 293355 379404 293421 379405
rect 293355 379340 293356 379404
rect 293420 379340 293421 379404
rect 293355 379339 293421 379340
rect 295931 379404 295997 379405
rect 295931 379340 295932 379404
rect 295996 379340 295997 379404
rect 295931 379339 295997 379340
rect 298507 379404 298573 379405
rect 298507 379340 298508 379404
rect 298572 379340 298573 379404
rect 298507 379339 298573 379340
rect 300899 379404 300965 379405
rect 300899 379340 300900 379404
rect 300964 379340 300965 379404
rect 300899 379339 300965 379340
rect 303475 379404 303541 379405
rect 303475 379340 303476 379404
rect 303540 379340 303541 379404
rect 303475 379339 303541 379340
rect 305867 379404 305933 379405
rect 305867 379340 305868 379404
rect 305932 379340 305933 379404
rect 305867 379339 305933 379340
rect 278451 379268 278517 379269
rect 278451 379204 278452 379268
rect 278516 379204 278517 379268
rect 278451 379203 278517 379204
rect 279187 379268 279253 379269
rect 279187 379204 279188 379268
rect 279252 379204 279253 379268
rect 279187 379203 279253 379204
rect 280843 379268 280909 379269
rect 280843 379204 280844 379268
rect 280908 379204 280909 379268
rect 280843 379203 280909 379204
rect 283419 379268 283485 379269
rect 283419 379204 283420 379268
rect 283484 379204 283485 379268
rect 283419 379203 283485 379204
rect 273483 378588 273549 378589
rect 273483 378524 273484 378588
rect 273548 378524 273549 378588
rect 273483 378523 273549 378524
rect 271794 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 272414 364394
rect 271794 364074 272414 364158
rect 271794 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 272414 364074
rect 271794 359308 272414 363838
rect 275514 368114 276134 379000
rect 275514 367878 275546 368114
rect 275782 367878 275866 368114
rect 276102 367878 276134 368114
rect 275514 367794 276134 367878
rect 275514 367558 275546 367794
rect 275782 367558 275866 367794
rect 276102 367558 276134 367794
rect 275514 359308 276134 367558
rect 279234 369954 279854 379000
rect 279234 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 279854 369954
rect 279234 369634 279854 369718
rect 279234 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 279854 369634
rect 279234 359308 279854 369398
rect 282954 373674 283574 379000
rect 282954 373438 282986 373674
rect 283222 373438 283306 373674
rect 283542 373438 283574 373674
rect 282954 373354 283574 373438
rect 282954 373118 282986 373354
rect 283222 373118 283306 373354
rect 283542 373118 283574 373354
rect 282954 359308 283574 373118
rect 289794 363454 290414 379000
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 359308 290414 362898
rect 293514 367174 294134 379000
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 359308 294134 366618
rect 297234 370894 297854 379000
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 359308 297854 370338
rect 300954 374614 301574 379000
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 359308 301574 374058
rect 307794 364394 308414 379000
rect 308630 378181 308690 380430
rect 311022 379405 311082 380430
rect 313414 380430 313500 380490
rect 315806 380430 315948 380490
rect 318382 380430 318532 380490
rect 320920 380490 320980 381106
rect 323368 380490 323428 381106
rect 325952 380490 326012 381106
rect 343224 380490 343284 381106
rect 320920 380430 321018 380490
rect 313414 379405 313474 380430
rect 315806 379405 315866 380430
rect 318382 379405 318442 380430
rect 311019 379404 311085 379405
rect 311019 379340 311020 379404
rect 311084 379340 311085 379404
rect 311019 379339 311085 379340
rect 313411 379404 313477 379405
rect 313411 379340 313412 379404
rect 313476 379340 313477 379404
rect 313411 379339 313477 379340
rect 315803 379404 315869 379405
rect 315803 379340 315804 379404
rect 315868 379340 315869 379404
rect 315803 379339 315869 379340
rect 318379 379404 318445 379405
rect 318379 379340 318380 379404
rect 318444 379340 318445 379404
rect 318379 379339 318445 379340
rect 308627 378180 308693 378181
rect 308627 378116 308628 378180
rect 308692 378116 308693 378180
rect 308627 378115 308693 378116
rect 307794 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 308414 364394
rect 307794 364074 308414 364158
rect 307794 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 308414 364074
rect 307794 359308 308414 363838
rect 311514 368114 312134 379000
rect 311514 367878 311546 368114
rect 311782 367878 311866 368114
rect 312102 367878 312134 368114
rect 311514 367794 312134 367878
rect 311514 367558 311546 367794
rect 311782 367558 311866 367794
rect 312102 367558 312134 367794
rect 311514 359308 312134 367558
rect 315234 369954 315854 379000
rect 315234 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 315854 369954
rect 315234 369634 315854 369718
rect 315234 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 315854 369634
rect 315234 359308 315854 369398
rect 318954 373674 319574 379000
rect 320958 378589 321018 380430
rect 323350 380430 323428 380490
rect 325926 380430 326012 380490
rect 343222 380430 343284 380490
rect 343360 380490 343420 381106
rect 343360 380430 343466 380490
rect 323350 379405 323410 380430
rect 325926 379405 325986 380430
rect 323347 379404 323413 379405
rect 323347 379340 323348 379404
rect 323412 379340 323413 379404
rect 323347 379339 323413 379340
rect 325923 379404 325989 379405
rect 325923 379340 325924 379404
rect 325988 379340 325989 379404
rect 325923 379339 325989 379340
rect 320955 378588 321021 378589
rect 320955 378524 320956 378588
rect 321020 378524 321021 378588
rect 320955 378523 321021 378524
rect 318954 373438 318986 373674
rect 319222 373438 319306 373674
rect 319542 373438 319574 373674
rect 318954 373354 319574 373438
rect 318954 373118 318986 373354
rect 319222 373118 319306 373354
rect 319542 373118 319574 373354
rect 318954 359308 319574 373118
rect 325794 363454 326414 379000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 359308 326414 362898
rect 329514 367174 330134 379000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 359308 330134 366618
rect 333234 370894 333854 379000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 359308 333854 370338
rect 336954 374614 337574 379000
rect 343222 378453 343282 380430
rect 343406 379405 343466 380430
rect 343403 379404 343469 379405
rect 343403 379340 343404 379404
rect 343468 379340 343469 379404
rect 343403 379339 343469 379340
rect 343219 378452 343285 378453
rect 343219 378388 343220 378452
rect 343284 378388 343285 378452
rect 343219 378387 343285 378388
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 359308 337574 374058
rect 343794 364394 344414 379000
rect 343794 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 344414 364394
rect 343794 364074 344414 364158
rect 343794 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 344414 364074
rect 343794 359308 344414 363838
rect 347514 368114 348134 379000
rect 347514 367878 347546 368114
rect 347782 367878 347866 368114
rect 348102 367878 348134 368114
rect 347514 367794 348134 367878
rect 347514 367558 347546 367794
rect 347782 367558 347866 367794
rect 348102 367558 348134 367794
rect 347514 359308 348134 367558
rect 351234 369954 351854 379000
rect 351234 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 351854 369954
rect 351234 369634 351854 369718
rect 351234 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 351854 369634
rect 351234 359308 351854 369398
rect 354954 373674 355574 379000
rect 354954 373438 354986 373674
rect 355222 373438 355306 373674
rect 355542 373438 355574 373674
rect 354954 373354 355574 373438
rect 354954 373118 354986 373354
rect 355222 373118 355306 373354
rect 355542 373118 355574 373354
rect 354954 359308 355574 373118
rect 338435 358868 338501 358869
rect 338435 358804 338436 358868
rect 338500 358804 338501 358868
rect 338435 358803 338501 358804
rect 339723 358868 339789 358869
rect 339723 358804 339724 358868
rect 339788 358804 339789 358868
rect 339723 358803 339789 358804
rect 350947 358868 351013 358869
rect 350947 358804 350948 358868
rect 351012 358804 351013 358868
rect 350947 358803 351013 358804
rect 338438 358050 338498 358803
rect 339726 358050 339786 358803
rect 350950 358050 351010 358803
rect 338438 357990 338524 358050
rect 338464 357202 338524 357990
rect 339688 357990 339786 358050
rect 350840 357990 351010 358050
rect 339688 357202 339748 357990
rect 350840 357202 350900 357990
rect 220272 345454 220620 345486
rect 220272 345218 220328 345454
rect 220564 345218 220620 345454
rect 220272 345134 220620 345218
rect 220272 344898 220328 345134
rect 220564 344898 220620 345134
rect 220272 344866 220620 344898
rect 356000 345454 356348 345486
rect 356000 345218 356056 345454
rect 356292 345218 356348 345454
rect 356000 345134 356348 345218
rect 356000 344898 356056 345134
rect 356292 344898 356348 345134
rect 356000 344866 356348 344898
rect 220952 327454 221300 327486
rect 220952 327218 221008 327454
rect 221244 327218 221300 327454
rect 220952 327134 221300 327218
rect 220952 326898 221008 327134
rect 221244 326898 221300 327134
rect 220952 326866 221300 326898
rect 355320 327454 355668 327486
rect 355320 327218 355376 327454
rect 355612 327218 355668 327454
rect 355320 327134 355668 327218
rect 355320 326898 355376 327134
rect 355612 326898 355668 327134
rect 355320 326866 355668 326898
rect 220272 309454 220620 309486
rect 220272 309218 220328 309454
rect 220564 309218 220620 309454
rect 220272 309134 220620 309218
rect 220272 308898 220328 309134
rect 220564 308898 220620 309134
rect 220272 308866 220620 308898
rect 356000 309454 356348 309486
rect 356000 309218 356056 309454
rect 356292 309218 356348 309454
rect 356000 309134 356348 309218
rect 356000 308898 356056 309134
rect 356292 308898 356348 309134
rect 356000 308866 356348 308898
rect 220952 291454 221300 291486
rect 220952 291218 221008 291454
rect 221244 291218 221300 291454
rect 220952 291134 221300 291218
rect 220952 290898 221008 291134
rect 221244 290898 221300 291134
rect 220952 290866 221300 290898
rect 355320 291454 355668 291486
rect 355320 291218 355376 291454
rect 355612 291218 355668 291454
rect 355320 291134 355668 291218
rect 355320 290898 355376 291134
rect 355612 290898 355668 291134
rect 355320 290866 355668 290898
rect 236056 273730 236116 274040
rect 237144 273730 237204 274040
rect 238232 273730 238292 274040
rect 239592 273730 239652 274040
rect 236056 273670 236562 273730
rect 221514 259174 222134 272000
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 252308 222134 258618
rect 225234 262894 225854 272000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 252308 225854 262338
rect 228954 266614 229574 272000
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 252308 229574 266058
rect 235794 256394 236414 272000
rect 236502 271421 236562 273670
rect 237054 273670 237204 273730
rect 238158 273670 238292 273730
rect 239262 273670 239652 273730
rect 240544 273730 240604 274040
rect 241768 273730 241828 274040
rect 243128 273730 243188 274040
rect 240544 273670 240610 273730
rect 236499 271420 236565 271421
rect 236499 271356 236500 271420
rect 236564 271356 236565 271420
rect 236499 271355 236565 271356
rect 237054 270605 237114 273670
rect 238158 270605 238218 273670
rect 237051 270604 237117 270605
rect 237051 270540 237052 270604
rect 237116 270540 237117 270604
rect 237051 270539 237117 270540
rect 238155 270604 238221 270605
rect 238155 270540 238156 270604
rect 238220 270540 238221 270604
rect 238155 270539 238221 270540
rect 239262 269789 239322 273670
rect 239259 269788 239325 269789
rect 239259 269724 239260 269788
rect 239324 269724 239325 269788
rect 239259 269723 239325 269724
rect 235794 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 236414 256394
rect 235794 256074 236414 256158
rect 235794 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 236414 256074
rect 235794 252308 236414 255838
rect 239514 260114 240134 272000
rect 240550 270197 240610 273670
rect 241654 273670 241828 273730
rect 242942 273670 243188 273730
rect 244216 273730 244276 274040
rect 245440 273730 245500 274040
rect 246528 273730 246588 274040
rect 244216 273670 244290 273730
rect 241654 270333 241714 273670
rect 242942 270605 243002 273670
rect 242939 270604 243005 270605
rect 242939 270540 242940 270604
rect 243004 270540 243005 270604
rect 242939 270539 243005 270540
rect 241651 270332 241717 270333
rect 241651 270268 241652 270332
rect 241716 270268 241717 270332
rect 241651 270267 241717 270268
rect 240547 270196 240613 270197
rect 240547 270132 240548 270196
rect 240612 270132 240613 270196
rect 240547 270131 240613 270132
rect 239514 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 240134 260114
rect 239514 259794 240134 259878
rect 239514 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 240134 259794
rect 239514 252308 240134 259558
rect 243234 261954 243854 272000
rect 244230 270741 244290 273670
rect 245334 273670 245500 273730
rect 246438 273670 246588 273730
rect 247616 273730 247676 274040
rect 248296 273730 248356 274040
rect 248704 273730 248764 274040
rect 247616 273670 247786 273730
rect 244227 270740 244293 270741
rect 244227 270676 244228 270740
rect 244292 270676 244293 270740
rect 244227 270675 244293 270676
rect 245334 270605 245394 273670
rect 246438 270605 246498 273670
rect 245331 270604 245397 270605
rect 245331 270540 245332 270604
rect 245396 270540 245397 270604
rect 245331 270539 245397 270540
rect 246435 270604 246501 270605
rect 246435 270540 246436 270604
rect 246500 270540 246501 270604
rect 246435 270539 246501 270540
rect 243234 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 243854 261954
rect 243234 261634 243854 261718
rect 243234 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 243854 261634
rect 243234 252308 243854 261398
rect 246954 265674 247574 272000
rect 247726 270605 247786 273670
rect 248278 273670 248356 273730
rect 248646 273670 248764 273730
rect 250064 273730 250124 274040
rect 250744 273730 250804 274040
rect 251288 273730 251348 274040
rect 252376 273730 252436 274040
rect 253464 273730 253524 274040
rect 250064 273670 250178 273730
rect 248278 271149 248338 273670
rect 248275 271148 248341 271149
rect 248275 271084 248276 271148
rect 248340 271084 248341 271148
rect 248275 271083 248341 271084
rect 248646 270605 248706 273670
rect 250118 270605 250178 273670
rect 250670 273670 250804 273730
rect 251222 273670 251348 273730
rect 252326 273670 252436 273730
rect 253430 273670 253524 273730
rect 253600 273730 253660 274040
rect 254552 273730 254612 274040
rect 255912 273730 255972 274040
rect 253600 273670 253674 273730
rect 250670 273325 250730 273670
rect 250667 273324 250733 273325
rect 250667 273260 250668 273324
rect 250732 273260 250733 273324
rect 250667 273259 250733 273260
rect 251222 270741 251282 273670
rect 251219 270740 251285 270741
rect 251219 270676 251220 270740
rect 251284 270676 251285 270740
rect 251219 270675 251285 270676
rect 252326 270605 252386 273670
rect 253430 270605 253490 273670
rect 253614 271149 253674 273670
rect 254534 273670 254612 273730
rect 255822 273670 255972 273730
rect 256048 273730 256108 274040
rect 257000 273730 257060 274040
rect 256048 273670 256250 273730
rect 253611 271148 253677 271149
rect 253611 271084 253612 271148
rect 253676 271084 253677 271148
rect 253611 271083 253677 271084
rect 247723 270604 247789 270605
rect 247723 270540 247724 270604
rect 247788 270540 247789 270604
rect 247723 270539 247789 270540
rect 248643 270604 248709 270605
rect 248643 270540 248644 270604
rect 248708 270540 248709 270604
rect 248643 270539 248709 270540
rect 250115 270604 250181 270605
rect 250115 270540 250116 270604
rect 250180 270540 250181 270604
rect 250115 270539 250181 270540
rect 252323 270604 252389 270605
rect 252323 270540 252324 270604
rect 252388 270540 252389 270604
rect 252323 270539 252389 270540
rect 253427 270604 253493 270605
rect 253427 270540 253428 270604
rect 253492 270540 253493 270604
rect 253427 270539 253493 270540
rect 246954 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 247574 265674
rect 246954 265354 247574 265438
rect 246954 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 247574 265354
rect 246954 252308 247574 265118
rect 253794 255454 254414 272000
rect 254534 270877 254594 273670
rect 254531 270876 254597 270877
rect 254531 270812 254532 270876
rect 254596 270812 254597 270876
rect 254531 270811 254597 270812
rect 255822 270741 255882 273670
rect 256190 271149 256250 273670
rect 256926 273670 257060 273730
rect 258088 273730 258148 274040
rect 258496 273730 258556 274040
rect 258088 273670 258274 273730
rect 256187 271148 256253 271149
rect 256187 271084 256188 271148
rect 256252 271084 256253 271148
rect 256187 271083 256253 271084
rect 255819 270740 255885 270741
rect 255819 270676 255820 270740
rect 255884 270676 255885 270740
rect 255819 270675 255885 270676
rect 256926 270605 256986 273670
rect 256923 270604 256989 270605
rect 256923 270540 256924 270604
rect 256988 270540 256989 270604
rect 256923 270539 256989 270540
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 252308 254414 254898
rect 257514 259174 258134 272000
rect 258214 271010 258274 273670
rect 258398 273670 258556 273730
rect 259448 273730 259508 274040
rect 260672 273730 260732 274040
rect 261080 273730 261140 274040
rect 259448 273670 259562 273730
rect 258398 271285 258458 273670
rect 258395 271284 258461 271285
rect 258395 271220 258396 271284
rect 258460 271220 258461 271284
rect 258395 271219 258461 271220
rect 258214 270950 258458 271010
rect 258398 270605 258458 270950
rect 259502 270605 259562 273670
rect 260606 273670 260732 273730
rect 260974 273670 261140 273730
rect 261760 273730 261820 274040
rect 262848 273730 262908 274040
rect 261760 273670 262138 273730
rect 260606 270741 260666 273670
rect 260974 271421 261034 273670
rect 260971 271420 261037 271421
rect 260971 271356 260972 271420
rect 261036 271356 261037 271420
rect 260971 271355 261037 271356
rect 260603 270740 260669 270741
rect 260603 270676 260604 270740
rect 260668 270676 260669 270740
rect 260603 270675 260669 270676
rect 258395 270604 258461 270605
rect 258395 270540 258396 270604
rect 258460 270540 258461 270604
rect 258395 270539 258461 270540
rect 259499 270604 259565 270605
rect 259499 270540 259500 270604
rect 259564 270540 259565 270604
rect 259499 270539 259565 270540
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 252308 258134 258618
rect 261234 262894 261854 272000
rect 262078 270605 262138 273670
rect 262814 273670 262908 273730
rect 263528 273730 263588 274040
rect 263936 273730 263996 274040
rect 265296 273730 265356 274040
rect 265976 273730 266036 274040
rect 263528 273670 263610 273730
rect 262814 270605 262874 273670
rect 263550 271829 263610 273670
rect 263918 273670 263996 273730
rect 265206 273670 265356 273730
rect 265942 273670 266036 273730
rect 263547 271828 263613 271829
rect 263547 271764 263548 271828
rect 263612 271764 263613 271828
rect 263547 271763 263613 271764
rect 263918 270605 263978 273670
rect 265206 272237 265266 273670
rect 265203 272236 265269 272237
rect 265203 272172 265204 272236
rect 265268 272172 265269 272236
rect 265203 272171 265269 272172
rect 262075 270604 262141 270605
rect 262075 270540 262076 270604
rect 262140 270540 262141 270604
rect 262075 270539 262141 270540
rect 262811 270604 262877 270605
rect 262811 270540 262812 270604
rect 262876 270540 262877 270604
rect 262811 270539 262877 270540
rect 263915 270604 263981 270605
rect 263915 270540 263916 270604
rect 263980 270540 263981 270604
rect 263915 270539 263981 270540
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 252308 261854 262338
rect 264954 266614 265574 272000
rect 265942 271285 266002 273670
rect 266384 273597 266444 274040
rect 267608 273730 267668 274040
rect 267598 273670 267668 273730
rect 268288 273730 268348 274040
rect 268696 273730 268756 274040
rect 268288 273670 268394 273730
rect 268696 273670 268762 273730
rect 266381 273596 266447 273597
rect 266381 273532 266382 273596
rect 266446 273532 266447 273596
rect 266381 273531 266447 273532
rect 265939 271284 266005 271285
rect 265939 271220 265940 271284
rect 266004 271220 266005 271284
rect 265939 271219 266005 271220
rect 267598 270605 267658 273670
rect 268334 271421 268394 273670
rect 268331 271420 268397 271421
rect 268331 271356 268332 271420
rect 268396 271356 268397 271420
rect 268331 271355 268397 271356
rect 268702 270605 268762 273670
rect 269784 273597 269844 274040
rect 271008 273730 271068 274040
rect 270910 273670 271068 273730
rect 269781 273596 269847 273597
rect 269781 273532 269782 273596
rect 269846 273532 269847 273596
rect 269781 273531 269847 273532
rect 270910 271829 270970 273670
rect 271144 273597 271204 274040
rect 272232 273730 272292 274040
rect 273320 273730 273380 274040
rect 273592 273730 273652 274040
rect 274408 273869 274468 274040
rect 274405 273868 274471 273869
rect 274405 273804 274406 273868
rect 274470 273804 274471 273868
rect 274405 273803 274471 273804
rect 275768 273730 275828 274040
rect 272232 273670 272626 273730
rect 271141 273596 271207 273597
rect 271141 273532 271142 273596
rect 271206 273532 271207 273596
rect 271141 273531 271207 273532
rect 270907 271828 270973 271829
rect 270907 271764 270908 271828
rect 270972 271764 270973 271828
rect 270907 271763 270973 271764
rect 267595 270604 267661 270605
rect 267595 270540 267596 270604
rect 267660 270540 267661 270604
rect 267595 270539 267661 270540
rect 268699 270604 268765 270605
rect 268699 270540 268700 270604
rect 268764 270540 268765 270604
rect 268699 270539 268765 270540
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 252308 265574 266058
rect 271794 256394 272414 272000
rect 272566 271829 272626 273670
rect 273302 273670 273380 273730
rect 273486 273670 273652 273730
rect 275326 273670 275828 273730
rect 276040 273730 276100 274040
rect 276992 273730 277052 274040
rect 276040 273670 276306 273730
rect 273302 273461 273362 273670
rect 273299 273460 273365 273461
rect 273299 273396 273300 273460
rect 273364 273396 273365 273460
rect 273299 273395 273365 273396
rect 272563 271828 272629 271829
rect 272563 271764 272564 271828
rect 272628 271764 272629 271828
rect 272563 271763 272629 271764
rect 273486 271557 273546 273670
rect 273483 271556 273549 271557
rect 273483 271492 273484 271556
rect 273548 271492 273549 271556
rect 273483 271491 273549 271492
rect 275326 271285 275386 273670
rect 275323 271284 275389 271285
rect 275323 271220 275324 271284
rect 275388 271220 275389 271284
rect 275323 271219 275389 271220
rect 271794 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 272414 256394
rect 271794 256074 272414 256158
rect 271794 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 272414 256074
rect 271794 252308 272414 255838
rect 275514 260114 276134 272000
rect 276246 271557 276306 273670
rect 276982 273670 277052 273730
rect 278080 273730 278140 274040
rect 278488 273730 278548 274040
rect 279168 273730 279228 274040
rect 280936 273730 280996 274040
rect 278080 273670 278146 273730
rect 276982 271829 277042 273670
rect 276979 271828 277045 271829
rect 276979 271764 276980 271828
rect 277044 271764 277045 271828
rect 276979 271763 277045 271764
rect 276243 271556 276309 271557
rect 276243 271492 276244 271556
rect 276308 271492 276309 271556
rect 276243 271491 276309 271492
rect 278086 271285 278146 273670
rect 278454 273670 278548 273730
rect 279006 273670 279228 273730
rect 280846 273670 280996 273730
rect 278454 271829 278514 273670
rect 278451 271828 278517 271829
rect 278451 271764 278452 271828
rect 278516 271764 278517 271828
rect 278451 271763 278517 271764
rect 278083 271284 278149 271285
rect 278083 271220 278084 271284
rect 278148 271220 278149 271284
rect 278083 271219 278149 271220
rect 279006 270877 279066 273670
rect 279003 270876 279069 270877
rect 279003 270812 279004 270876
rect 279068 270812 279069 270876
rect 279003 270811 279069 270812
rect 275514 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 276134 260114
rect 275514 259794 276134 259878
rect 275514 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 276134 259794
rect 275514 252308 276134 259558
rect 279234 261954 279854 272000
rect 280846 271829 280906 273670
rect 283520 273597 283580 274040
rect 285968 273730 286028 274040
rect 288280 273730 288340 274040
rect 291000 273730 291060 274040
rect 293448 273730 293508 274040
rect 285968 273670 286058 273730
rect 283517 273596 283583 273597
rect 283517 273532 283518 273596
rect 283582 273532 283583 273596
rect 283517 273531 283583 273532
rect 285998 272917 286058 273670
rect 288206 273670 288340 273730
rect 290966 273670 291060 273730
rect 293358 273670 293508 273730
rect 295896 273730 295956 274040
rect 298480 273730 298540 274040
rect 300928 273730 300988 274040
rect 303512 273730 303572 274040
rect 305960 273730 306020 274040
rect 295896 273670 295994 273730
rect 298480 273670 298570 273730
rect 288206 272917 288266 273670
rect 290966 272917 291026 273670
rect 293358 272917 293418 273670
rect 295934 272917 295994 273670
rect 298510 273053 298570 273670
rect 300902 273670 300988 273730
rect 303478 273670 303572 273730
rect 305870 273670 306020 273730
rect 308544 273730 308604 274040
rect 310992 273730 311052 274040
rect 313440 273730 313500 274040
rect 315888 273730 315948 274040
rect 318472 273730 318532 274040
rect 308544 273670 308690 273730
rect 310992 273670 311082 273730
rect 298507 273052 298573 273053
rect 298507 272988 298508 273052
rect 298572 272988 298573 273052
rect 298507 272987 298573 272988
rect 285995 272916 286061 272917
rect 285995 272852 285996 272916
rect 286060 272852 286061 272916
rect 285995 272851 286061 272852
rect 288203 272916 288269 272917
rect 288203 272852 288204 272916
rect 288268 272852 288269 272916
rect 288203 272851 288269 272852
rect 290963 272916 291029 272917
rect 290963 272852 290964 272916
rect 291028 272852 291029 272916
rect 290963 272851 291029 272852
rect 293355 272916 293421 272917
rect 293355 272852 293356 272916
rect 293420 272852 293421 272916
rect 293355 272851 293421 272852
rect 295931 272916 295997 272917
rect 295931 272852 295932 272916
rect 295996 272852 295997 272916
rect 295931 272851 295997 272852
rect 300902 272781 300962 273670
rect 303478 272781 303538 273670
rect 305870 272917 305930 273670
rect 305867 272916 305933 272917
rect 305867 272852 305868 272916
rect 305932 272852 305933 272916
rect 305867 272851 305933 272852
rect 300899 272780 300965 272781
rect 300899 272716 300900 272780
rect 300964 272716 300965 272780
rect 300899 272715 300965 272716
rect 303475 272780 303541 272781
rect 303475 272716 303476 272780
rect 303540 272716 303541 272780
rect 303475 272715 303541 272716
rect 280843 271828 280909 271829
rect 280843 271764 280844 271828
rect 280908 271764 280909 271828
rect 280843 271763 280909 271764
rect 279234 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 279854 261954
rect 279234 261634 279854 261718
rect 279234 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 279854 261634
rect 279234 252308 279854 261398
rect 282954 265674 283574 272000
rect 282954 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 283574 265674
rect 282954 265354 283574 265438
rect 282954 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 283574 265354
rect 282954 252308 283574 265118
rect 289794 255454 290414 272000
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 252308 290414 254898
rect 293514 259174 294134 272000
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 252308 294134 258618
rect 297234 262894 297854 272000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 252308 297854 262338
rect 300954 266614 301574 272000
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 252308 301574 266058
rect 307794 256394 308414 272000
rect 308630 271829 308690 273670
rect 311022 272645 311082 273670
rect 313414 273670 313500 273730
rect 315070 273670 315948 273730
rect 318382 273670 318532 273730
rect 320920 273730 320980 274040
rect 323368 273730 323428 274040
rect 325952 273730 326012 274040
rect 343224 273730 343284 274040
rect 320920 273670 321018 273730
rect 311019 272644 311085 272645
rect 311019 272580 311020 272644
rect 311084 272580 311085 272644
rect 311019 272579 311085 272580
rect 308627 271828 308693 271829
rect 308627 271764 308628 271828
rect 308692 271764 308693 271828
rect 308627 271763 308693 271764
rect 307794 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 308414 256394
rect 307794 256074 308414 256158
rect 307794 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 308414 256074
rect 307794 252308 308414 255838
rect 311514 260114 312134 272000
rect 313414 271149 313474 273670
rect 315070 271693 315130 273670
rect 318382 273189 318442 273670
rect 318379 273188 318445 273189
rect 318379 273124 318380 273188
rect 318444 273124 318445 273188
rect 318379 273123 318445 273124
rect 320958 272645 321018 273670
rect 323350 273670 323428 273730
rect 325742 273670 326012 273730
rect 343222 273670 343284 273730
rect 343360 273730 343420 274040
rect 343360 273670 343466 273730
rect 320955 272644 321021 272645
rect 320955 272580 320956 272644
rect 321020 272580 321021 272644
rect 320955 272579 321021 272580
rect 315067 271692 315133 271693
rect 315067 271628 315068 271692
rect 315132 271628 315133 271692
rect 315067 271627 315133 271628
rect 313411 271148 313477 271149
rect 313411 271084 313412 271148
rect 313476 271084 313477 271148
rect 313411 271083 313477 271084
rect 311514 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 312134 260114
rect 311514 259794 312134 259878
rect 311514 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 312134 259794
rect 311514 252308 312134 259558
rect 315234 261954 315854 272000
rect 315234 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 315854 261954
rect 315234 261634 315854 261718
rect 315234 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 315854 261634
rect 315234 252308 315854 261398
rect 318954 265674 319574 272000
rect 323350 270469 323410 273670
rect 325742 272370 325802 273670
rect 325558 272310 325802 272370
rect 325558 271013 325618 272310
rect 325555 271012 325621 271013
rect 325555 270948 325556 271012
rect 325620 270948 325621 271012
rect 325555 270947 325621 270948
rect 323347 270468 323413 270469
rect 323347 270404 323348 270468
rect 323412 270404 323413 270468
rect 323347 270403 323413 270404
rect 318954 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 319574 265674
rect 318954 265354 319574 265438
rect 318954 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 319574 265354
rect 318954 252308 319574 265118
rect 325794 255454 326414 272000
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 252308 326414 254898
rect 329514 259174 330134 272000
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 252308 330134 258618
rect 333234 262894 333854 272000
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 252308 333854 262338
rect 336954 266614 337574 272000
rect 343222 271421 343282 273670
rect 343406 271829 343466 273670
rect 343403 271828 343469 271829
rect 343403 271764 343404 271828
rect 343468 271764 343469 271828
rect 343403 271763 343469 271764
rect 343219 271420 343285 271421
rect 343219 271356 343220 271420
rect 343284 271356 343285 271420
rect 343219 271355 343285 271356
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 252308 337574 266058
rect 343794 256394 344414 272000
rect 343794 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 344414 256394
rect 343794 256074 344414 256158
rect 343794 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 344414 256074
rect 339723 253468 339789 253469
rect 339723 253404 339724 253468
rect 339788 253404 339789 253468
rect 339723 253403 339789 253404
rect 338435 253060 338501 253061
rect 338435 252996 338436 253060
rect 338500 252996 338501 253060
rect 338435 252995 338501 252996
rect 338438 250610 338498 252995
rect 339726 250610 339786 253403
rect 343794 252308 344414 255838
rect 347514 260114 348134 272000
rect 347514 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 348134 260114
rect 347514 259794 348134 259878
rect 347514 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 348134 259794
rect 347514 252308 348134 259558
rect 351234 261954 351854 272000
rect 351234 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 351854 261954
rect 351234 261634 351854 261718
rect 351234 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 351854 261634
rect 350947 253196 351013 253197
rect 350947 253132 350948 253196
rect 351012 253132 351013 253196
rect 350947 253131 351013 253132
rect 350950 250610 351010 253131
rect 351234 252308 351854 261398
rect 354954 265674 355574 272000
rect 354954 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 355574 265674
rect 354954 265354 355574 265438
rect 354954 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 355574 265354
rect 354954 252308 355574 265118
rect 338438 250550 338524 250610
rect 338464 250240 338524 250550
rect 339688 250550 339786 250610
rect 350840 250550 351010 250610
rect 339688 250240 339748 250550
rect 350840 250240 350900 250550
rect 220272 237454 220620 237486
rect 220272 237218 220328 237454
rect 220564 237218 220620 237454
rect 220272 237134 220620 237218
rect 220272 236898 220328 237134
rect 220564 236898 220620 237134
rect 220272 236866 220620 236898
rect 356000 237454 356348 237486
rect 356000 237218 356056 237454
rect 356292 237218 356348 237454
rect 356000 237134 356348 237218
rect 356000 236898 356056 237134
rect 356292 236898 356348 237134
rect 356000 236866 356348 236898
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 201454 220620 201486
rect 220272 201218 220328 201454
rect 220564 201218 220620 201454
rect 220272 201134 220620 201218
rect 220272 200898 220328 201134
rect 220564 200898 220620 201134
rect 220272 200866 220620 200898
rect 356000 201454 356348 201486
rect 356000 201218 356056 201454
rect 356292 201218 356348 201454
rect 356000 201134 356348 201218
rect 356000 200898 356056 201134
rect 356292 200898 356348 201134
rect 356000 200866 356348 200898
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 166290 236116 167106
rect 237144 166290 237204 167106
rect 238232 166290 238292 167106
rect 236056 166230 236194 166290
rect 236134 165613 236194 166230
rect 237054 166230 237204 166290
rect 238158 166230 238292 166290
rect 239592 166290 239652 167106
rect 240544 166290 240604 167106
rect 241768 166290 241828 167106
rect 243128 166290 243188 167106
rect 244216 167010 244276 167106
rect 245440 167010 245500 167106
rect 246528 167010 246588 167106
rect 247616 167010 247676 167106
rect 248296 167010 248356 167106
rect 248704 167010 248764 167106
rect 244216 166950 244474 167010
rect 244216 166910 244290 166950
rect 239592 166230 239690 166290
rect 240544 166230 240610 166290
rect 236131 165612 236197 165613
rect 236131 165548 236132 165612
rect 236196 165548 236197 165612
rect 236131 165547 236197 165548
rect 221514 151174 222134 165000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 145308 222134 150618
rect 225234 154894 225854 165000
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 145308 225854 154338
rect 228954 158614 229574 165000
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 145308 229574 158058
rect 235794 148394 236414 165000
rect 237054 164253 237114 166230
rect 238158 164253 238218 166230
rect 239630 165613 239690 166230
rect 239627 165612 239693 165613
rect 239627 165548 239628 165612
rect 239692 165548 239693 165612
rect 239627 165547 239693 165548
rect 237051 164252 237117 164253
rect 237051 164188 237052 164252
rect 237116 164188 237117 164252
rect 237051 164187 237117 164188
rect 238155 164252 238221 164253
rect 238155 164188 238156 164252
rect 238220 164188 238221 164252
rect 238155 164187 238221 164188
rect 235794 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 236414 148394
rect 235794 148074 236414 148158
rect 235794 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 236414 148074
rect 235794 145308 236414 147838
rect 239514 152114 240134 165000
rect 240550 164253 240610 166230
rect 241654 166230 241828 166290
rect 243126 166230 243188 166290
rect 241654 164253 241714 166230
rect 243126 165613 243186 166230
rect 243123 165612 243189 165613
rect 243123 165548 243124 165612
rect 243188 165548 243189 165612
rect 243123 165547 243189 165548
rect 240547 164252 240613 164253
rect 240547 164188 240548 164252
rect 240612 164188 240613 164252
rect 240547 164187 240613 164188
rect 241651 164252 241717 164253
rect 241651 164188 241652 164252
rect 241716 164188 241717 164252
rect 241651 164187 241717 164188
rect 239514 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 240134 152114
rect 239514 151794 240134 151878
rect 239514 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 240134 151794
rect 239514 145308 240134 151558
rect 243234 155834 243854 165000
rect 244414 164389 244474 166950
rect 245334 166950 245500 167010
rect 246438 166950 246588 167010
rect 247542 166950 247676 167010
rect 248278 166950 248356 167010
rect 248646 166950 248764 167010
rect 250064 167010 250124 167106
rect 250744 167010 250804 167106
rect 251288 167010 251348 167106
rect 252376 167010 252436 167106
rect 253464 167010 253524 167106
rect 250064 166950 250178 167010
rect 244411 164388 244477 164389
rect 244411 164324 244412 164388
rect 244476 164324 244477 164388
rect 244411 164323 244477 164324
rect 245334 164253 245394 166950
rect 246438 164253 246498 166950
rect 247542 165613 247602 166950
rect 247539 165612 247605 165613
rect 247539 165548 247540 165612
rect 247604 165548 247605 165612
rect 247539 165547 247605 165548
rect 245331 164252 245397 164253
rect 245331 164188 245332 164252
rect 245396 164188 245397 164252
rect 245331 164187 245397 164188
rect 246435 164252 246501 164253
rect 246435 164188 246436 164252
rect 246500 164188 246501 164252
rect 246435 164187 246501 164188
rect 243234 155598 243266 155834
rect 243502 155598 243586 155834
rect 243822 155598 243854 155834
rect 243234 155514 243854 155598
rect 243234 155278 243266 155514
rect 243502 155278 243586 155514
rect 243822 155278 243854 155514
rect 243234 145308 243854 155278
rect 246954 157674 247574 165000
rect 248278 164933 248338 166950
rect 248275 164932 248341 164933
rect 248275 164868 248276 164932
rect 248340 164868 248341 164932
rect 248275 164867 248341 164868
rect 248646 164253 248706 166950
rect 250118 164253 250178 166950
rect 250670 166950 250804 167010
rect 251222 166950 251348 167010
rect 252326 166950 252436 167010
rect 253430 166950 253524 167010
rect 253600 167010 253660 167106
rect 254552 167010 254612 167106
rect 255912 167010 255972 167106
rect 253600 166950 253674 167010
rect 250670 164933 250730 166950
rect 250667 164932 250733 164933
rect 250667 164868 250668 164932
rect 250732 164868 250733 164932
rect 250667 164867 250733 164868
rect 251222 164253 251282 166950
rect 252326 164389 252386 166950
rect 252323 164388 252389 164389
rect 252323 164324 252324 164388
rect 252388 164324 252389 164388
rect 252323 164323 252389 164324
rect 253430 164253 253490 166950
rect 253614 164933 253674 166950
rect 254534 166950 254612 167010
rect 255822 166950 255972 167010
rect 256048 167010 256108 167106
rect 257000 167010 257060 167106
rect 258088 167010 258148 167106
rect 258496 167010 258556 167106
rect 256048 166950 256250 167010
rect 253611 164932 253677 164933
rect 253611 164868 253612 164932
rect 253676 164868 253677 164932
rect 253611 164867 253677 164868
rect 248643 164252 248709 164253
rect 248643 164188 248644 164252
rect 248708 164188 248709 164252
rect 248643 164187 248709 164188
rect 250115 164252 250181 164253
rect 250115 164188 250116 164252
rect 250180 164188 250181 164252
rect 250115 164187 250181 164188
rect 251219 164252 251285 164253
rect 251219 164188 251220 164252
rect 251284 164188 251285 164252
rect 251219 164187 251285 164188
rect 253427 164252 253493 164253
rect 253427 164188 253428 164252
rect 253492 164188 253493 164252
rect 253427 164187 253493 164188
rect 246954 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 247574 157674
rect 246954 157354 247574 157438
rect 246954 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 247574 157354
rect 246954 145308 247574 157118
rect 253794 147454 254414 165000
rect 254534 164253 254594 166950
rect 255822 164253 255882 166950
rect 256190 165613 256250 166950
rect 256926 166950 257060 167010
rect 258030 166950 258148 167010
rect 258398 166950 258556 167010
rect 259448 167010 259508 167106
rect 260672 167010 260732 167106
rect 261080 167010 261140 167106
rect 261760 167010 261820 167106
rect 262848 167010 262908 167106
rect 259448 166950 259562 167010
rect 256187 165612 256253 165613
rect 256187 165548 256188 165612
rect 256252 165548 256253 165612
rect 256187 165547 256253 165548
rect 256926 164253 256986 166950
rect 258030 165613 258090 166950
rect 258027 165612 258093 165613
rect 258027 165548 258028 165612
rect 258092 165548 258093 165612
rect 258027 165547 258093 165548
rect 254531 164252 254597 164253
rect 254531 164188 254532 164252
rect 254596 164188 254597 164252
rect 254531 164187 254597 164188
rect 255819 164252 255885 164253
rect 255819 164188 255820 164252
rect 255884 164188 255885 164252
rect 255819 164187 255885 164188
rect 256923 164252 256989 164253
rect 256923 164188 256924 164252
rect 256988 164188 256989 164252
rect 256923 164187 256989 164188
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 145308 254414 146898
rect 257514 151174 258134 165000
rect 258398 164933 258458 166950
rect 258395 164932 258461 164933
rect 258395 164868 258396 164932
rect 258460 164868 258461 164932
rect 258395 164867 258461 164868
rect 259502 164253 259562 166950
rect 260606 166950 260732 167010
rect 260974 166950 261140 167010
rect 261710 166950 261820 167010
rect 262814 166950 262908 167010
rect 263528 167010 263588 167106
rect 263936 167010 263996 167106
rect 265296 167010 265356 167106
rect 265976 167010 266036 167106
rect 263528 166950 263794 167010
rect 260606 164389 260666 166950
rect 260974 166429 261034 166950
rect 260971 166428 261037 166429
rect 260971 166364 260972 166428
rect 261036 166364 261037 166428
rect 260971 166363 261037 166364
rect 261710 165613 261770 166950
rect 261707 165612 261773 165613
rect 261707 165548 261708 165612
rect 261772 165548 261773 165612
rect 261707 165547 261773 165548
rect 260603 164388 260669 164389
rect 260603 164324 260604 164388
rect 260668 164324 260669 164388
rect 260603 164323 260669 164324
rect 259499 164252 259565 164253
rect 259499 164188 259500 164252
rect 259564 164188 259565 164252
rect 259499 164187 259565 164188
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 145308 258134 150618
rect 261234 154894 261854 165000
rect 262814 164253 262874 166950
rect 263734 165205 263794 166950
rect 263918 166950 263996 167010
rect 265206 166950 265356 167010
rect 265942 166950 266036 167010
rect 266384 167010 266444 167106
rect 267608 167010 267668 167106
rect 266384 166950 266554 167010
rect 263731 165204 263797 165205
rect 263731 165140 263732 165204
rect 263796 165140 263797 165204
rect 263731 165139 263797 165140
rect 263918 164253 263978 166950
rect 265206 165205 265266 166950
rect 265942 166429 266002 166950
rect 265939 166428 266005 166429
rect 265939 166364 265940 166428
rect 266004 166364 266005 166428
rect 265939 166363 266005 166364
rect 265203 165204 265269 165205
rect 265203 165140 265204 165204
rect 265268 165140 265269 165204
rect 265203 165139 265269 165140
rect 262811 164252 262877 164253
rect 262811 164188 262812 164252
rect 262876 164188 262877 164252
rect 262811 164187 262877 164188
rect 263915 164252 263981 164253
rect 263915 164188 263916 164252
rect 263980 164188 263981 164252
rect 263915 164187 263981 164188
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 145308 261854 154338
rect 264954 158614 265574 165000
rect 266494 164389 266554 166950
rect 267598 166950 267668 167010
rect 268288 167010 268348 167106
rect 268696 167010 268756 167106
rect 269784 167010 269844 167106
rect 271008 167010 271068 167106
rect 268288 166950 268394 167010
rect 268696 166950 268762 167010
rect 269784 166950 269866 167010
rect 266491 164388 266557 164389
rect 266491 164324 266492 164388
rect 266556 164324 266557 164388
rect 266491 164323 266557 164324
rect 267598 164253 267658 166950
rect 268334 165205 268394 166950
rect 268331 165204 268397 165205
rect 268331 165140 268332 165204
rect 268396 165140 268397 165204
rect 268331 165139 268397 165140
rect 268702 164253 268762 166950
rect 269806 164253 269866 166950
rect 270910 166950 271068 167010
rect 271144 167010 271204 167106
rect 272232 167010 272292 167106
rect 273320 167010 273380 167106
rect 273592 167010 273652 167106
rect 274408 167010 274468 167106
rect 275768 167010 275828 167106
rect 271144 166950 271338 167010
rect 270910 166293 270970 166950
rect 270907 166292 270973 166293
rect 270907 166228 270908 166292
rect 270972 166228 270973 166292
rect 270907 166227 270973 166228
rect 271278 164253 271338 166950
rect 272198 166950 272292 167010
rect 273302 166950 273380 167010
rect 273486 166950 273652 167010
rect 274406 166950 274468 167010
rect 275694 166950 275828 167010
rect 276040 167010 276100 167106
rect 276992 167010 277052 167106
rect 276040 166950 276122 167010
rect 272198 165205 272258 166950
rect 272195 165204 272261 165205
rect 272195 165140 272196 165204
rect 272260 165140 272261 165204
rect 272195 165139 272261 165140
rect 267595 164252 267661 164253
rect 267595 164188 267596 164252
rect 267660 164188 267661 164252
rect 267595 164187 267661 164188
rect 268699 164252 268765 164253
rect 268699 164188 268700 164252
rect 268764 164188 268765 164252
rect 268699 164187 268765 164188
rect 269803 164252 269869 164253
rect 269803 164188 269804 164252
rect 269868 164188 269869 164252
rect 269803 164187 269869 164188
rect 271275 164252 271341 164253
rect 271275 164188 271276 164252
rect 271340 164188 271341 164252
rect 271275 164187 271341 164188
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 145308 265574 158058
rect 271794 148394 272414 165000
rect 273302 164253 273362 166950
rect 273486 165069 273546 166950
rect 273483 165068 273549 165069
rect 273483 165004 273484 165068
rect 273548 165004 273549 165068
rect 273483 165003 273549 165004
rect 274406 164389 274466 166950
rect 275694 165205 275754 166950
rect 276062 165205 276122 166950
rect 276982 166950 277052 167010
rect 278080 167010 278140 167106
rect 278488 167010 278548 167106
rect 278080 166950 278146 167010
rect 275691 165204 275757 165205
rect 275691 165140 275692 165204
rect 275756 165140 275757 165204
rect 275691 165139 275757 165140
rect 276059 165204 276125 165205
rect 276059 165140 276060 165204
rect 276124 165140 276125 165204
rect 276059 165139 276125 165140
rect 274403 164388 274469 164389
rect 274403 164324 274404 164388
rect 274468 164324 274469 164388
rect 274403 164323 274469 164324
rect 273299 164252 273365 164253
rect 273299 164188 273300 164252
rect 273364 164188 273365 164252
rect 273299 164187 273365 164188
rect 271794 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 272414 148394
rect 271794 148074 272414 148158
rect 271794 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 272414 148074
rect 271794 145308 272414 147838
rect 275514 152114 276134 165000
rect 276982 164253 277042 166950
rect 278086 164253 278146 166950
rect 278454 166950 278548 167010
rect 279168 167010 279228 167106
rect 280936 167010 280996 167106
rect 279168 166950 279250 167010
rect 278454 165613 278514 166950
rect 278451 165612 278517 165613
rect 278451 165548 278452 165612
rect 278516 165548 278517 165612
rect 278451 165547 278517 165548
rect 279190 165205 279250 166950
rect 280846 166950 280996 167010
rect 280846 165613 280906 166950
rect 283520 166290 283580 167106
rect 283422 166230 283580 166290
rect 285968 166293 286028 167106
rect 288280 166701 288340 167106
rect 291000 166701 291060 167106
rect 293448 167010 293508 167106
rect 293358 166950 293508 167010
rect 295896 167010 295956 167106
rect 298480 167010 298540 167106
rect 300928 167010 300988 167106
rect 295896 166950 295994 167010
rect 298480 166950 298570 167010
rect 288277 166700 288343 166701
rect 288277 166636 288278 166700
rect 288342 166636 288343 166700
rect 288277 166635 288343 166636
rect 290997 166700 291063 166701
rect 290997 166636 290998 166700
rect 291062 166636 291063 166700
rect 290997 166635 291063 166636
rect 293358 166429 293418 166950
rect 293355 166428 293421 166429
rect 293355 166364 293356 166428
rect 293420 166364 293421 166428
rect 293355 166363 293421 166364
rect 295934 166293 295994 166950
rect 298510 166429 298570 166950
rect 300902 166950 300988 167010
rect 298507 166428 298573 166429
rect 298507 166364 298508 166428
rect 298572 166364 298573 166428
rect 298507 166363 298573 166364
rect 285968 166292 286061 166293
rect 285968 166230 285996 166292
rect 283422 165613 283482 166230
rect 285995 166228 285996 166230
rect 286060 166228 286061 166292
rect 285995 166227 286061 166228
rect 295931 166292 295997 166293
rect 295931 166228 295932 166292
rect 295996 166228 295997 166292
rect 295931 166227 295997 166228
rect 300902 165613 300962 166950
rect 303512 166565 303572 167106
rect 305960 166837 306020 167106
rect 305957 166836 306023 166837
rect 305957 166772 305958 166836
rect 306022 166772 306023 166836
rect 308544 166834 308604 167106
rect 305957 166771 306023 166772
rect 308446 166774 308604 166834
rect 310992 166834 311052 167106
rect 313440 166837 313500 167106
rect 313437 166836 313503 166837
rect 310992 166774 311082 166834
rect 303509 166564 303575 166565
rect 303509 166500 303510 166564
rect 303574 166500 303575 166564
rect 303509 166499 303575 166500
rect 308446 165613 308506 166774
rect 280843 165612 280909 165613
rect 280843 165548 280844 165612
rect 280908 165548 280909 165612
rect 280843 165547 280909 165548
rect 283419 165612 283485 165613
rect 283419 165548 283420 165612
rect 283484 165548 283485 165612
rect 283419 165547 283485 165548
rect 300899 165612 300965 165613
rect 300899 165548 300900 165612
rect 300964 165548 300965 165612
rect 300899 165547 300965 165548
rect 308443 165612 308509 165613
rect 308443 165548 308444 165612
rect 308508 165548 308509 165612
rect 308443 165547 308509 165548
rect 311022 165341 311082 166774
rect 313437 166772 313438 166836
rect 313502 166772 313503 166836
rect 315888 166834 315948 167106
rect 318472 166834 318532 167106
rect 313437 166771 313503 166772
rect 315806 166774 315948 166834
rect 318382 166774 318532 166834
rect 320920 166834 320980 167106
rect 323368 166834 323428 167106
rect 320920 166774 321018 166834
rect 315806 165477 315866 166774
rect 315803 165476 315869 165477
rect 315803 165412 315804 165476
rect 315868 165412 315869 165476
rect 315803 165411 315869 165412
rect 311019 165340 311085 165341
rect 311019 165276 311020 165340
rect 311084 165276 311085 165340
rect 311019 165275 311085 165276
rect 279187 165204 279253 165205
rect 279187 165140 279188 165204
rect 279252 165140 279253 165204
rect 279187 165139 279253 165140
rect 276979 164252 277045 164253
rect 276979 164188 276980 164252
rect 277044 164188 277045 164252
rect 276979 164187 277045 164188
rect 278083 164252 278149 164253
rect 278083 164188 278084 164252
rect 278148 164188 278149 164252
rect 278083 164187 278149 164188
rect 275514 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 276134 152114
rect 275514 151794 276134 151878
rect 275514 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 276134 151794
rect 275514 145308 276134 151558
rect 279234 155834 279854 165000
rect 279234 155598 279266 155834
rect 279502 155598 279586 155834
rect 279822 155598 279854 155834
rect 279234 155514 279854 155598
rect 279234 155278 279266 155514
rect 279502 155278 279586 155514
rect 279822 155278 279854 155514
rect 279234 145308 279854 155278
rect 282954 157674 283574 165000
rect 282954 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 283574 157674
rect 282954 157354 283574 157438
rect 282954 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 283574 157354
rect 282954 145308 283574 157118
rect 289794 147454 290414 165000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 145308 290414 146898
rect 293514 151174 294134 165000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 145308 294134 150618
rect 297234 154894 297854 165000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 145308 297854 154338
rect 300954 158614 301574 165000
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 145308 301574 158058
rect 307794 148394 308414 165000
rect 307794 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 308414 148394
rect 307794 148074 308414 148158
rect 307794 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 308414 148074
rect 307794 145308 308414 147838
rect 311514 152114 312134 165000
rect 311514 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 312134 152114
rect 311514 151794 312134 151878
rect 311514 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 312134 151794
rect 311514 145308 312134 151558
rect 315234 155834 315854 165000
rect 318382 164253 318442 166774
rect 320958 165613 321018 166774
rect 323350 166774 323428 166834
rect 320955 165612 321021 165613
rect 320955 165548 320956 165612
rect 321020 165548 321021 165612
rect 320955 165547 321021 165548
rect 318379 164252 318445 164253
rect 318379 164188 318380 164252
rect 318444 164188 318445 164252
rect 318379 164187 318445 164188
rect 315234 155598 315266 155834
rect 315502 155598 315586 155834
rect 315822 155598 315854 155834
rect 315234 155514 315854 155598
rect 315234 155278 315266 155514
rect 315502 155278 315586 155514
rect 315822 155278 315854 155514
rect 315234 145308 315854 155278
rect 318954 157674 319574 165000
rect 323350 164797 323410 166774
rect 325952 166290 326012 167106
rect 343224 166290 343284 167106
rect 325926 166230 326012 166290
rect 343222 166230 343284 166290
rect 343360 166290 343420 167106
rect 356654 166973 356714 484875
rect 356651 166972 356717 166973
rect 356651 166908 356652 166972
rect 356716 166908 356717 166972
rect 356651 166907 356717 166908
rect 343360 166230 343466 166290
rect 325926 165613 325986 166230
rect 343222 165613 343282 166230
rect 343406 165613 343466 166230
rect 325923 165612 325989 165613
rect 325923 165548 325924 165612
rect 325988 165548 325989 165612
rect 325923 165547 325989 165548
rect 343219 165612 343285 165613
rect 343219 165548 343220 165612
rect 343284 165548 343285 165612
rect 343219 165547 343285 165548
rect 343403 165612 343469 165613
rect 343403 165548 343404 165612
rect 343468 165548 343469 165612
rect 343403 165547 343469 165548
rect 323347 164796 323413 164797
rect 323347 164732 323348 164796
rect 323412 164732 323413 164796
rect 323347 164731 323413 164732
rect 318954 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 319574 157674
rect 318954 157354 319574 157438
rect 318954 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 319574 157354
rect 318954 145308 319574 157118
rect 325794 147454 326414 165000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 145308 326414 146898
rect 329514 151174 330134 165000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 145308 330134 150618
rect 333234 154894 333854 165000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 145308 333854 154338
rect 336954 158614 337574 165000
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 145308 337574 158058
rect 343794 148394 344414 165000
rect 343794 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 344414 148394
rect 343794 148074 344414 148158
rect 343794 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 344414 148074
rect 343794 145308 344414 147838
rect 347514 152114 348134 165000
rect 347514 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 348134 152114
rect 347514 151794 348134 151878
rect 347514 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 348134 151794
rect 347514 145308 348134 151558
rect 351234 155834 351854 165000
rect 351234 155598 351266 155834
rect 351502 155598 351586 155834
rect 351822 155598 351854 155834
rect 351234 155514 351854 155598
rect 351234 155278 351266 155514
rect 351502 155278 351586 155514
rect 351822 155278 351854 155514
rect 351234 145308 351854 155278
rect 354954 157674 355574 165000
rect 354954 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 355574 157674
rect 354954 157354 355574 157438
rect 354954 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 355574 157354
rect 354954 145308 355574 157118
rect 338435 144940 338501 144941
rect 338435 144876 338436 144940
rect 338500 144876 338501 144940
rect 338435 144875 338501 144876
rect 339723 144940 339789 144941
rect 339723 144876 339724 144940
rect 339788 144876 339789 144940
rect 339723 144875 339789 144876
rect 350947 144940 351013 144941
rect 350947 144876 350948 144940
rect 351012 144876 351013 144940
rect 350947 144875 351013 144876
rect 338438 143850 338498 144875
rect 339726 143850 339786 144875
rect 350950 143850 351010 144875
rect 338438 143790 338524 143850
rect 338464 143202 338524 143790
rect 339688 143790 339786 143850
rect 350840 143790 351010 143850
rect 339688 143202 339748 143790
rect 350840 143202 350900 143790
rect 220272 129454 220620 129486
rect 220272 129218 220328 129454
rect 220564 129218 220620 129454
rect 220272 129134 220620 129218
rect 220272 128898 220328 129134
rect 220564 128898 220620 129134
rect 220272 128866 220620 128898
rect 356000 129454 356348 129486
rect 356000 129218 356056 129454
rect 356292 129218 356348 129454
rect 356000 129134 356348 129218
rect 356000 128898 356056 129134
rect 356292 128898 356348 129134
rect 356000 128866 356348 128898
rect 220952 111454 221300 111486
rect 220952 111218 221008 111454
rect 221244 111218 221300 111454
rect 220952 111134 221300 111218
rect 220952 110898 221008 111134
rect 221244 110898 221300 111134
rect 220952 110866 221300 110898
rect 355320 111454 355668 111486
rect 355320 111218 355376 111454
rect 355612 111218 355668 111454
rect 355320 111134 355668 111218
rect 355320 110898 355376 111134
rect 355612 110898 355668 111134
rect 355320 110866 355668 110898
rect 220272 93454 220620 93486
rect 220272 93218 220328 93454
rect 220564 93218 220620 93454
rect 220272 93134 220620 93218
rect 220272 92898 220328 93134
rect 220564 92898 220620 93134
rect 220272 92866 220620 92898
rect 356000 93454 356348 93486
rect 356000 93218 356056 93454
rect 356292 93218 356348 93454
rect 356000 93134 356348 93218
rect 356000 92898 356056 93134
rect 356292 92898 356348 93134
rect 356000 92866 356348 92898
rect 220952 75454 221300 75486
rect 220952 75218 221008 75454
rect 221244 75218 221300 75454
rect 220952 75134 221300 75218
rect 220952 74898 221008 75134
rect 221244 74898 221300 75134
rect 220952 74866 221300 74898
rect 355320 75454 355668 75486
rect 355320 75218 355376 75454
rect 355612 75218 355668 75454
rect 355320 75134 355668 75218
rect 355320 74898 355376 75134
rect 355612 74898 355668 75134
rect 355320 74866 355668 74898
rect 236056 59805 236116 60106
rect 237144 59805 237204 60106
rect 236053 59804 236119 59805
rect 236053 59740 236054 59804
rect 236118 59740 236119 59804
rect 236053 59739 236119 59740
rect 237141 59804 237207 59805
rect 237141 59740 237142 59804
rect 237206 59740 237207 59804
rect 237141 59739 237207 59740
rect 238232 59530 238292 60106
rect 239592 59530 239652 60106
rect 238158 59470 238292 59530
rect 239262 59470 239652 59530
rect 240544 59530 240604 60106
rect 241768 59530 241828 60106
rect 243128 59530 243188 60106
rect 240544 59470 240610 59530
rect 219939 56404 220005 56405
rect 219939 56340 219940 56404
rect 220004 56340 220005 56404
rect 219939 56339 220005 56340
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 238158 57901 238218 59470
rect 239262 57901 239322 59470
rect 238155 57900 238221 57901
rect 238155 57836 238156 57900
rect 238220 57836 238221 57900
rect 238155 57835 238221 57836
rect 239259 57900 239325 57901
rect 239259 57836 239260 57900
rect 239324 57836 239325 57900
rect 239259 57835 239325 57836
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 240550 57901 240610 59470
rect 241654 59470 241828 59530
rect 242942 59470 243188 59530
rect 244216 59530 244276 60106
rect 245440 59530 245500 60106
rect 246528 59530 246588 60106
rect 244216 59470 244290 59530
rect 241654 57901 241714 59470
rect 242942 57901 243002 59470
rect 240547 57900 240613 57901
rect 240547 57836 240548 57900
rect 240612 57836 240613 57900
rect 240547 57835 240613 57836
rect 241651 57900 241717 57901
rect 241651 57836 241652 57900
rect 241716 57836 241717 57900
rect 241651 57835 241717 57836
rect 242939 57900 243005 57901
rect 242939 57836 242940 57900
rect 243004 57836 243005 57900
rect 242939 57835 243005 57836
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 244230 57901 244290 59470
rect 245334 59470 245500 59530
rect 246438 59470 246588 59530
rect 247616 59530 247676 60106
rect 248296 59530 248356 60106
rect 248704 59530 248764 60106
rect 247616 59470 247786 59530
rect 245334 57901 245394 59470
rect 246438 57901 246498 59470
rect 244227 57900 244293 57901
rect 244227 57836 244228 57900
rect 244292 57836 244293 57900
rect 244227 57835 244293 57836
rect 245331 57900 245397 57901
rect 245331 57836 245332 57900
rect 245396 57836 245397 57900
rect 245331 57835 245397 57836
rect 246435 57900 246501 57901
rect 246435 57836 246436 57900
rect 246500 57836 246501 57900
rect 246435 57835 246501 57836
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 247726 57901 247786 59470
rect 248278 59470 248356 59530
rect 248646 59470 248764 59530
rect 250064 59530 250124 60106
rect 250744 59530 250804 60106
rect 251288 59530 251348 60106
rect 252376 59530 252436 60106
rect 253464 59530 253524 60106
rect 250064 59470 250178 59530
rect 247723 57900 247789 57901
rect 247723 57836 247724 57900
rect 247788 57836 247789 57900
rect 247723 57835 247789 57836
rect 248278 57221 248338 59470
rect 248646 57901 248706 59470
rect 250118 57901 250178 59470
rect 250670 59470 250804 59530
rect 251222 59470 251348 59530
rect 252326 59470 252436 59530
rect 253430 59470 253524 59530
rect 253600 59530 253660 60106
rect 254552 59530 254612 60106
rect 255912 59805 255972 60106
rect 255909 59804 255975 59805
rect 255909 59740 255910 59804
rect 255974 59740 255975 59804
rect 255909 59739 255975 59740
rect 256048 59530 256108 60106
rect 257000 59805 257060 60106
rect 256997 59804 257063 59805
rect 256997 59740 256998 59804
rect 257062 59740 257063 59804
rect 256997 59739 257063 59740
rect 258088 59530 258148 60106
rect 258496 59530 258556 60106
rect 253600 59470 253674 59530
rect 250670 58581 250730 59470
rect 250667 58580 250733 58581
rect 250667 58516 250668 58580
rect 250732 58516 250733 58580
rect 250667 58515 250733 58516
rect 248643 57900 248709 57901
rect 248643 57836 248644 57900
rect 248708 57836 248709 57900
rect 248643 57835 248709 57836
rect 250115 57900 250181 57901
rect 250115 57836 250116 57900
rect 250180 57836 250181 57900
rect 250115 57835 250181 57836
rect 251222 57493 251282 59470
rect 252326 57493 252386 59470
rect 253430 57493 253490 59470
rect 253614 58717 253674 59470
rect 254534 59470 254612 59530
rect 256006 59470 256108 59530
rect 257846 59470 258148 59530
rect 258398 59470 258556 59530
rect 259448 59530 259508 60106
rect 260672 59669 260732 60106
rect 260669 59668 260735 59669
rect 260669 59604 260670 59668
rect 260734 59604 260735 59668
rect 260669 59603 260735 59604
rect 261080 59530 261140 60106
rect 261760 59530 261820 60106
rect 262848 59805 262908 60106
rect 262845 59804 262911 59805
rect 262845 59740 262846 59804
rect 262910 59740 262911 59804
rect 262845 59739 262911 59740
rect 259448 59470 259562 59530
rect 253611 58716 253677 58717
rect 253611 58652 253612 58716
rect 253676 58652 253677 58716
rect 253611 58651 253677 58652
rect 251219 57492 251285 57493
rect 251219 57428 251220 57492
rect 251284 57428 251285 57492
rect 251219 57427 251285 57428
rect 252323 57492 252389 57493
rect 252323 57428 252324 57492
rect 252388 57428 252389 57492
rect 252323 57427 252389 57428
rect 253427 57492 253493 57493
rect 253427 57428 253428 57492
rect 253492 57428 253493 57492
rect 253427 57427 253493 57428
rect 248275 57220 248341 57221
rect 248275 57156 248276 57220
rect 248340 57156 248341 57220
rect 248275 57155 248341 57156
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 254534 57493 254594 59470
rect 256006 57901 256066 59470
rect 257846 58445 257906 59470
rect 257843 58444 257909 58445
rect 257843 58380 257844 58444
rect 257908 58380 257909 58444
rect 257843 58379 257909 58380
rect 256003 57900 256069 57901
rect 256003 57836 256004 57900
rect 256068 57836 256069 57900
rect 256003 57835 256069 57836
rect 254531 57492 254597 57493
rect 254531 57428 254532 57492
rect 254596 57428 254597 57492
rect 254531 57427 254597 57428
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 258398 57765 258458 59470
rect 259502 59397 259562 59470
rect 260974 59470 261140 59530
rect 261710 59470 261820 59530
rect 263528 59533 263588 60106
rect 263528 59532 263613 59533
rect 263528 59470 263548 59532
rect 259499 59396 259565 59397
rect 259499 59332 259500 59396
rect 259564 59332 259565 59396
rect 259499 59331 259565 59332
rect 258395 57764 258461 57765
rect 258395 57700 258396 57764
rect 258460 57700 258461 57764
rect 258395 57699 258461 57700
rect 260974 57085 261034 59470
rect 261710 59397 261770 59470
rect 263547 59468 263548 59470
rect 263612 59468 263613 59532
rect 263936 59530 263996 60106
rect 265296 59530 265356 60106
rect 265976 59530 266036 60106
rect 266384 59530 266444 60106
rect 267608 59530 267668 60106
rect 263547 59467 263613 59468
rect 263918 59470 263996 59530
rect 265206 59470 265356 59530
rect 265942 59470 266036 59530
rect 266310 59470 266444 59530
rect 267598 59470 267668 59530
rect 268288 59530 268348 60106
rect 268696 59530 268756 60106
rect 269784 59530 269844 60106
rect 271008 59666 271068 60106
rect 270910 59606 271068 59666
rect 268288 59470 268394 59530
rect 268696 59470 268762 59530
rect 269784 59470 269866 59530
rect 261707 59396 261773 59397
rect 261707 59332 261708 59396
rect 261772 59332 261773 59396
rect 261707 59331 261773 59332
rect 260971 57084 261037 57085
rect 260971 57020 260972 57084
rect 261036 57020 261037 57084
rect 260971 57019 261037 57020
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 263918 57765 263978 59470
rect 265206 58173 265266 59470
rect 265203 58172 265269 58173
rect 265203 58108 265204 58172
rect 265268 58108 265269 58172
rect 265203 58107 265269 58108
rect 263915 57764 263981 57765
rect 263915 57700 263916 57764
rect 263980 57700 263981 57764
rect 263915 57699 263981 57700
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 265942 57357 266002 59470
rect 266310 57493 266370 59470
rect 267598 57765 267658 59470
rect 268334 58853 268394 59470
rect 268331 58852 268397 58853
rect 268331 58788 268332 58852
rect 268396 58788 268397 58852
rect 268331 58787 268397 58788
rect 268702 57765 268762 59470
rect 269806 57765 269866 59470
rect 270910 57901 270970 59606
rect 271144 59530 271204 60106
rect 272232 59530 272292 60106
rect 273320 59530 273380 60106
rect 273592 59666 273652 60106
rect 271094 59470 271204 59530
rect 272198 59470 272292 59530
rect 273302 59470 273380 59530
rect 273486 59606 273652 59666
rect 271094 57901 271154 59470
rect 272198 58173 272258 59470
rect 272195 58172 272261 58173
rect 272195 58108 272196 58172
rect 272260 58108 272261 58172
rect 272195 58107 272261 58108
rect 270907 57900 270973 57901
rect 270907 57836 270908 57900
rect 270972 57836 270973 57900
rect 270907 57835 270973 57836
rect 271091 57900 271157 57901
rect 271091 57836 271092 57900
rect 271156 57836 271157 57900
rect 271091 57835 271157 57836
rect 267595 57764 267661 57765
rect 267595 57700 267596 57764
rect 267660 57700 267661 57764
rect 267595 57699 267661 57700
rect 268699 57764 268765 57765
rect 268699 57700 268700 57764
rect 268764 57700 268765 57764
rect 268699 57699 268765 57700
rect 269803 57764 269869 57765
rect 269803 57700 269804 57764
rect 269868 57700 269869 57764
rect 269803 57699 269869 57700
rect 266307 57492 266373 57493
rect 266307 57428 266308 57492
rect 266372 57428 266373 57492
rect 266307 57427 266373 57428
rect 271794 57454 272414 58000
rect 273302 57901 273362 59470
rect 273299 57900 273365 57901
rect 273299 57836 273300 57900
rect 273364 57836 273365 57900
rect 273299 57835 273365 57836
rect 265939 57356 266005 57357
rect 265939 57292 265940 57356
rect 266004 57292 266005 57356
rect 265939 57291 266005 57292
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 273486 56269 273546 59606
rect 274408 59530 274468 60106
rect 275768 59666 275828 60106
rect 274406 59470 274468 59530
rect 275694 59606 275828 59666
rect 276040 59666 276100 60106
rect 276040 59606 276122 59666
rect 274406 57765 274466 59470
rect 275694 58173 275754 59606
rect 276062 59261 276122 59606
rect 276992 59530 277052 60106
rect 278080 59530 278140 60106
rect 278488 59530 278548 60106
rect 276982 59470 277052 59530
rect 277902 59470 278140 59530
rect 278454 59470 278548 59530
rect 279168 59530 279228 60106
rect 280936 59530 280996 60106
rect 279168 59470 279250 59530
rect 276059 59260 276125 59261
rect 276059 59196 276060 59260
rect 276124 59196 276125 59260
rect 276059 59195 276125 59196
rect 275691 58172 275757 58173
rect 275691 58108 275692 58172
rect 275756 58108 275757 58172
rect 275691 58107 275757 58108
rect 274403 57764 274469 57765
rect 274403 57700 274404 57764
rect 274468 57700 274469 57764
rect 274403 57699 274469 57700
rect 273483 56268 273549 56269
rect 273483 56204 273484 56268
rect 273548 56204 273549 56268
rect 273483 56203 273549 56204
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 276982 57901 277042 59470
rect 277902 57990 277962 59470
rect 277166 57930 277962 57990
rect 276979 57900 277045 57901
rect 276979 57836 276980 57900
rect 277044 57836 277045 57900
rect 276979 57835 277045 57836
rect 277166 56133 277226 57930
rect 278454 57629 278514 59470
rect 279190 59261 279250 59470
rect 280846 59470 280996 59530
rect 283520 59530 283580 60106
rect 285968 59530 286028 60106
rect 288280 59530 288340 60106
rect 291000 59530 291060 60106
rect 293448 59530 293508 60106
rect 283520 59470 283850 59530
rect 285968 59470 286058 59530
rect 279187 59260 279253 59261
rect 279187 59196 279188 59260
rect 279252 59196 279253 59260
rect 279187 59195 279253 59196
rect 280846 59125 280906 59470
rect 280843 59124 280909 59125
rect 280843 59060 280844 59124
rect 280908 59060 280909 59124
rect 280843 59059 280909 59060
rect 278451 57628 278517 57629
rect 278451 57564 278452 57628
rect 278516 57564 278517 57628
rect 278451 57563 278517 57564
rect 277163 56132 277229 56133
rect 277163 56068 277164 56132
rect 277228 56068 277229 56132
rect 277163 56067 277229 56068
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 283790 56677 283850 59470
rect 285998 58989 286058 59470
rect 288206 59470 288340 59530
rect 290966 59470 291060 59530
rect 293358 59470 293508 59530
rect 295896 59530 295956 60106
rect 298480 59530 298540 60106
rect 300928 59530 300988 60106
rect 303512 59530 303572 60106
rect 305960 59530 306020 60106
rect 308544 59669 308604 60106
rect 308541 59668 308607 59669
rect 308541 59604 308542 59668
rect 308606 59604 308607 59668
rect 308541 59603 308607 59604
rect 295896 59470 295994 59530
rect 298480 59470 298570 59530
rect 285995 58988 286061 58989
rect 285995 58924 285996 58988
rect 286060 58924 286061 58988
rect 285995 58923 286061 58924
rect 288206 57901 288266 59470
rect 290966 59261 291026 59470
rect 290963 59260 291029 59261
rect 290963 59196 290964 59260
rect 291028 59196 291029 59260
rect 290963 59195 291029 59196
rect 288203 57900 288269 57901
rect 288203 57836 288204 57900
rect 288268 57836 288269 57900
rect 288203 57835 288269 57836
rect 283787 56676 283853 56677
rect 283787 56612 283788 56676
rect 283852 56612 283853 56676
rect 283787 56611 283853 56612
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 293358 57901 293418 59470
rect 293355 57900 293421 57901
rect 293355 57836 293356 57900
rect 293420 57836 293421 57900
rect 293355 57835 293421 57836
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 295934 57901 295994 59470
rect 295931 57900 295997 57901
rect 295931 57836 295932 57900
rect 295996 57836 295997 57900
rect 295931 57835 295997 57836
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 298510 57901 298570 59470
rect 300902 59470 300988 59530
rect 303478 59470 303572 59530
rect 305870 59470 306020 59530
rect 310992 59530 311052 60106
rect 313440 59530 313500 60106
rect 315888 59669 315948 60106
rect 315885 59668 315951 59669
rect 315885 59604 315886 59668
rect 315950 59604 315951 59668
rect 318472 59666 318532 60106
rect 315885 59603 315951 59604
rect 318382 59606 318532 59666
rect 310992 59470 311082 59530
rect 300902 59261 300962 59470
rect 300899 59260 300965 59261
rect 300899 59196 300900 59260
rect 300964 59196 300965 59260
rect 300899 59195 300965 59196
rect 298507 57900 298573 57901
rect 298507 57836 298508 57900
rect 298572 57836 298573 57900
rect 298507 57835 298573 57836
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 303478 57901 303538 59470
rect 305870 57901 305930 59470
rect 303475 57900 303541 57901
rect 303475 57836 303476 57900
rect 303540 57836 303541 57900
rect 303475 57835 303541 57836
rect 305867 57900 305933 57901
rect 305867 57836 305868 57900
rect 305932 57836 305933 57900
rect 305867 57835 305933 57836
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 311022 57901 311082 59470
rect 313414 59470 313500 59530
rect 311019 57900 311085 57901
rect 311019 57836 311020 57900
rect 311084 57836 311085 57900
rect 311019 57835 311085 57836
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 313414 57901 313474 59470
rect 313411 57900 313477 57901
rect 313411 57836 313412 57900
rect 313476 57836 313477 57900
rect 313411 57835 313477 57836
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 318382 57901 318442 59606
rect 320920 59530 320980 60106
rect 323368 59530 323428 60106
rect 325952 59530 326012 60106
rect 343224 59530 343284 60106
rect 320920 59470 321018 59530
rect 320958 59261 321018 59470
rect 323350 59470 323428 59530
rect 325926 59470 326012 59530
rect 343222 59470 343284 59530
rect 343360 59530 343420 60106
rect 343360 59470 343466 59530
rect 320955 59260 321021 59261
rect 320955 59196 320956 59260
rect 321020 59196 321021 59260
rect 320955 59195 321021 59196
rect 318379 57900 318445 57901
rect 318379 57836 318380 57900
rect 318444 57836 318445 57900
rect 318379 57835 318445 57836
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 323350 57901 323410 59470
rect 325926 59261 325986 59470
rect 325923 59260 325989 59261
rect 325923 59196 325924 59260
rect 325988 59196 325989 59260
rect 325923 59195 325989 59196
rect 323347 57900 323413 57901
rect 323347 57836 323348 57900
rect 323412 57836 323413 57900
rect 323347 57835 323413 57836
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 343222 57901 343282 59470
rect 343406 57901 343466 59470
rect 357942 59261 358002 485691
rect 360699 483716 360765 483717
rect 360699 483652 360700 483716
rect 360764 483652 360765 483716
rect 360699 483651 360765 483652
rect 359411 475420 359477 475421
rect 359411 475356 359412 475420
rect 359476 475356 359477 475420
rect 359411 475355 359477 475356
rect 358123 474468 358189 474469
rect 358123 474404 358124 474468
rect 358188 474404 358189 474468
rect 358123 474403 358189 474404
rect 357939 59260 358005 59261
rect 357939 59196 357940 59260
rect 358004 59196 358005 59260
rect 357939 59195 358005 59196
rect 343219 57900 343285 57901
rect 343219 57836 343220 57900
rect 343284 57836 343285 57900
rect 343219 57835 343285 57836
rect 343403 57900 343469 57901
rect 343403 57836 343404 57900
rect 343468 57836 343469 57900
rect 343403 57835 343469 57836
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 358126 57765 358186 474403
rect 359414 273325 359474 475355
rect 359779 474604 359845 474605
rect 359779 474540 359780 474604
rect 359844 474540 359845 474604
rect 359779 474539 359845 474540
rect 359595 468484 359661 468485
rect 359595 468420 359596 468484
rect 359660 468420 359661 468484
rect 359595 468419 359661 468420
rect 359411 273324 359477 273325
rect 359411 273260 359412 273324
rect 359476 273260 359477 273324
rect 359411 273259 359477 273260
rect 359598 273189 359658 468419
rect 359782 378045 359842 474539
rect 359963 467124 360029 467125
rect 359963 467060 359964 467124
rect 360028 467060 360029 467124
rect 359963 467059 360029 467060
rect 359966 381581 360026 467059
rect 359963 381580 360029 381581
rect 359963 381516 359964 381580
rect 360028 381516 360029 381580
rect 359963 381515 360029 381516
rect 359779 378044 359845 378045
rect 359779 377980 359780 378044
rect 359844 377980 359845 378044
rect 359779 377979 359845 377980
rect 359595 273188 359661 273189
rect 359595 273124 359596 273188
rect 359660 273124 359661 273188
rect 359595 273123 359661 273124
rect 358123 57764 358189 57765
rect 358123 57700 358124 57764
rect 358188 57700 358189 57764
rect 358123 57699 358189 57700
rect 360702 56677 360762 483651
rect 360886 149157 360946 516699
rect 361794 507454 362414 520000
rect 363459 515404 363525 515405
rect 363459 515340 363460 515404
rect 363524 515340 363525 515404
rect 363459 515339 363525 515340
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 360883 149156 360949 149157
rect 360883 149092 360884 149156
rect 360948 149092 360949 149156
rect 360883 149091 360949 149092
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 360699 56676 360765 56677
rect 360699 56612 360700 56676
rect 360764 56612 360765 56676
rect 360699 56611 360765 56612
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 363462 3773 363522 515339
rect 365514 511174 366134 520000
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 363643 491876 363709 491877
rect 363643 491812 363644 491876
rect 363708 491812 363709 491876
rect 363643 491811 363709 491812
rect 363459 3772 363525 3773
rect 363459 3708 363460 3772
rect 363524 3708 363525 3772
rect 363459 3707 363525 3708
rect 363646 3501 363706 491811
rect 364931 485620 364997 485621
rect 364931 485556 364932 485620
rect 364996 485556 364997 485620
rect 364931 485555 364997 485556
rect 364379 479636 364445 479637
rect 364379 479572 364380 479636
rect 364444 479572 364445 479636
rect 364379 479571 364445 479572
rect 364382 379541 364442 479571
rect 364379 379540 364445 379541
rect 364379 379476 364380 379540
rect 364444 379476 364445 379540
rect 364379 379475 364445 379476
rect 364934 58853 364994 485555
rect 365514 475174 366134 510618
rect 369234 514894 369854 520000
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 367691 490516 367757 490517
rect 367691 490452 367692 490516
rect 367756 490452 367757 490516
rect 367691 490451 367757 490452
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 364931 58852 364997 58853
rect 364931 58788 364932 58852
rect 364996 58788 364997 58852
rect 364931 58787 364997 58788
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 363643 3500 363709 3501
rect 363643 3436 363644 3500
rect 363708 3436 363709 3500
rect 363643 3435 363709 3436
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 -2266 366134 6618
rect 367694 3365 367754 490451
rect 367875 487796 367941 487797
rect 367875 487732 367876 487796
rect 367940 487732 367941 487796
rect 367875 487731 367941 487732
rect 367878 3637 367938 487731
rect 369234 478894 369854 514338
rect 372954 518614 373574 520000
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 371739 485484 371805 485485
rect 371739 485420 371740 485484
rect 371804 485420 371805 485484
rect 371739 485419 371805 485420
rect 370083 480860 370149 480861
rect 370083 480796 370084 480860
rect 370148 480796 370149 480860
rect 370083 480795 370149 480796
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 370086 376821 370146 480795
rect 370451 476916 370517 476917
rect 370451 476852 370452 476916
rect 370516 476852 370517 476916
rect 370451 476851 370517 476852
rect 370083 376820 370149 376821
rect 370083 376756 370084 376820
rect 370148 376756 370149 376820
rect 370083 376755 370149 376756
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 370454 57493 370514 476851
rect 371742 58989 371802 485419
rect 372954 482614 373574 518058
rect 379794 489454 380414 520000
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 373763 485348 373829 485349
rect 373763 485284 373764 485348
rect 373828 485284 373829 485348
rect 373763 485283 373829 485284
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 371739 58988 371805 58989
rect 371739 58924 371740 58988
rect 371804 58924 371805 58988
rect 371739 58923 371805 58924
rect 370451 57492 370517 57493
rect 370451 57428 370452 57492
rect 370516 57428 370517 57492
rect 370451 57427 370517 57428
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 367875 3636 367941 3637
rect 367875 3572 367876 3636
rect 367940 3572 367941 3636
rect 367875 3571 367941 3572
rect 367691 3364 367757 3365
rect 367691 3300 367692 3364
rect 367756 3300 367757 3364
rect 367691 3299 367757 3300
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 86058
rect 373766 59125 373826 485283
rect 374499 485212 374565 485213
rect 374499 485148 374500 485212
rect 374564 485148 374565 485212
rect 374499 485147 374565 485148
rect 373763 59124 373829 59125
rect 373763 59060 373764 59124
rect 373828 59060 373829 59124
rect 373763 59059 373829 59060
rect 374502 58717 374562 485147
rect 375971 485076 376037 485077
rect 375971 485012 375972 485076
rect 376036 485012 376037 485076
rect 375971 485011 376037 485012
rect 375419 482492 375485 482493
rect 375419 482428 375420 482492
rect 375484 482428 375485 482492
rect 375419 482427 375485 482428
rect 374867 480996 374933 480997
rect 374867 480932 374868 480996
rect 374932 480932 374933 480996
rect 374867 480931 374933 480932
rect 374683 474196 374749 474197
rect 374683 474132 374684 474196
rect 374748 474132 374749 474196
rect 374683 474131 374749 474132
rect 374499 58716 374565 58717
rect 374499 58652 374500 58716
rect 374564 58652 374565 58716
rect 374499 58651 374565 58652
rect 374686 57629 374746 474131
rect 374870 165205 374930 480931
rect 375422 375189 375482 482427
rect 375419 375188 375485 375189
rect 375419 375124 375420 375188
rect 375484 375124 375485 375188
rect 375419 375123 375485 375124
rect 374867 165204 374933 165205
rect 374867 165140 374868 165204
rect 374932 165140 374933 165204
rect 374867 165139 374933 165140
rect 375974 58581 376034 485011
rect 377443 483988 377509 483989
rect 377443 483924 377444 483988
rect 377508 483924 377509 483988
rect 377443 483923 377509 483924
rect 377259 483852 377325 483853
rect 377259 483788 377260 483852
rect 377324 483788 377325 483852
rect 377259 483787 377325 483788
rect 376155 482356 376221 482357
rect 376155 482292 376156 482356
rect 376220 482292 376221 482356
rect 376155 482291 376221 482292
rect 376158 68101 376218 482291
rect 376891 477052 376957 477053
rect 376891 476988 376892 477052
rect 376956 476988 376957 477052
rect 376891 476987 376957 476988
rect 376894 378997 376954 476987
rect 376891 378996 376957 378997
rect 376891 378932 376892 378996
rect 376956 378932 376957 378996
rect 376891 378931 376957 378932
rect 376894 378181 376954 378931
rect 376891 378180 376957 378181
rect 376891 378116 376892 378180
rect 376956 378116 376957 378180
rect 376891 378115 376957 378116
rect 377262 271421 377322 483787
rect 377446 376685 377506 483923
rect 378731 478276 378797 478277
rect 378731 478212 378732 478276
rect 378796 478212 378797 478276
rect 378731 478211 378797 478212
rect 378179 476780 378245 476781
rect 378179 476716 378180 476780
rect 378244 476716 378245 476780
rect 378179 476715 378245 476716
rect 377627 475556 377693 475557
rect 377627 475492 377628 475556
rect 377692 475492 377693 475556
rect 377627 475491 377693 475492
rect 377630 382397 377690 475491
rect 377627 382396 377693 382397
rect 377627 382332 377628 382396
rect 377692 382332 377693 382396
rect 377627 382331 377693 382332
rect 377443 376684 377509 376685
rect 377443 376620 377444 376684
rect 377508 376620 377509 376684
rect 377443 376619 377509 376620
rect 377443 375324 377509 375325
rect 377443 375260 377444 375324
rect 377508 375260 377509 375324
rect 377443 375259 377509 375260
rect 377446 273461 377506 375259
rect 377995 374780 378061 374781
rect 377995 374716 377996 374780
rect 378060 374716 378061 374780
rect 377995 374715 378061 374716
rect 377443 273460 377509 273461
rect 377443 273396 377444 273460
rect 377508 273396 377509 273460
rect 377443 273395 377509 273396
rect 377811 273460 377877 273461
rect 377811 273396 377812 273460
rect 377876 273396 377877 273460
rect 377811 273395 377877 273396
rect 377814 273053 377874 273395
rect 377811 273052 377877 273053
rect 377811 272988 377812 273052
rect 377876 272988 377877 273052
rect 377811 272987 377877 272988
rect 377259 271420 377325 271421
rect 377259 271356 377260 271420
rect 377324 271356 377325 271420
rect 377259 271355 377325 271356
rect 377998 265029 378058 374715
rect 378182 273461 378242 476715
rect 378179 273460 378245 273461
rect 378179 273396 378180 273460
rect 378244 273396 378245 273460
rect 378179 273395 378245 273396
rect 377995 265028 378061 265029
rect 377995 264964 377996 265028
rect 378060 264964 378061 265028
rect 377995 264963 378061 264964
rect 377995 252516 378061 252517
rect 377995 252452 377996 252516
rect 378060 252452 378061 252516
rect 377995 252451 378061 252452
rect 377627 148340 377693 148341
rect 377627 148276 377628 148340
rect 377692 148276 377693 148340
rect 377627 148275 377693 148276
rect 376155 68100 376221 68101
rect 376155 68036 376156 68100
rect 376220 68036 376221 68100
rect 376155 68035 376221 68036
rect 375971 58580 376037 58581
rect 375971 58516 375972 58580
rect 376036 58516 376037 58580
rect 375971 58515 376037 58516
rect 374683 57628 374749 57629
rect 374683 57564 374684 57628
rect 374748 57564 374749 57628
rect 374683 57563 374749 57564
rect 377630 56269 377690 148275
rect 377998 146301 378058 252451
rect 377995 146300 378061 146301
rect 377995 146236 377996 146300
rect 378060 146236 378061 146300
rect 377995 146235 378061 146236
rect 377811 145756 377877 145757
rect 377811 145692 377812 145756
rect 377876 145692 377877 145756
rect 377811 145691 377877 145692
rect 377627 56268 377693 56269
rect 377627 56204 377628 56268
rect 377692 56204 377693 56268
rect 377627 56203 377693 56204
rect 377814 55997 377874 145691
rect 378734 57085 378794 478211
rect 379467 474332 379533 474333
rect 379467 474268 379468 474332
rect 379532 474330 379533 474332
rect 379532 474270 379714 474330
rect 379532 474268 379533 474270
rect 379467 474267 379533 474268
rect 378915 474060 378981 474061
rect 378915 473996 378916 474060
rect 378980 473996 378981 474060
rect 378915 473995 378981 473996
rect 378918 57221 378978 473995
rect 379099 472564 379165 472565
rect 379099 472500 379100 472564
rect 379164 472500 379165 472564
rect 379099 472499 379165 472500
rect 379102 57357 379162 472499
rect 379654 171150 379714 474270
rect 379794 466308 380414 488898
rect 383514 493174 384134 520000
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 466308 384134 492618
rect 387234 496894 387854 520000
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 466308 387854 496338
rect 390954 500614 391574 520000
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 466308 391574 500058
rect 397794 507454 398414 520000
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 466308 398414 470898
rect 401514 511174 402134 520000
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 466308 402134 474618
rect 405234 514894 405854 520000
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 466308 405854 478338
rect 408954 518614 409574 520000
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 466308 409574 482058
rect 415794 489454 416414 520000
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 466308 416414 488898
rect 419514 493174 420134 520000
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 466308 420134 492618
rect 423234 496894 423854 520000
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 466308 423854 496338
rect 426954 500614 427574 520000
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 466308 427574 500058
rect 433794 507454 434414 520000
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 466308 434414 470898
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 466308 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 466308 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 466308 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 466308 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 630000 459854 640338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 630000 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 630000 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 630000 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 630000 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 630000 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 630000 488414 632898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 630000 492134 636618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 630000 495854 640338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 630000 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 630000 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 630000 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 476067 627876 476133 627877
rect 476067 627812 476068 627876
rect 476132 627812 476133 627876
rect 476067 627811 476133 627812
rect 488579 627876 488645 627877
rect 488579 627812 488580 627876
rect 488644 627812 488645 627876
rect 488579 627811 488645 627812
rect 506611 627876 506677 627877
rect 506611 627812 506612 627876
rect 506676 627812 506677 627876
rect 506611 627811 506677 627812
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 466308 456134 492618
rect 459234 568894 459854 576000
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 466308 459854 496338
rect 462954 572614 463574 576000
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 466308 463574 500058
rect 469794 543454 470414 576000
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 466308 470414 470898
rect 473514 547174 474134 576000
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 476070 491877 476130 627811
rect 479568 597454 479888 597486
rect 479568 597218 479610 597454
rect 479846 597218 479888 597454
rect 479568 597134 479888 597218
rect 479568 596898 479610 597134
rect 479846 596898 479888 597134
rect 479568 596866 479888 596898
rect 477234 550894 477854 576000
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 476067 491876 476133 491877
rect 476067 491812 476068 491876
rect 476132 491812 476133 491876
rect 476067 491811 476133 491812
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 466308 474134 474618
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 466308 477854 478338
rect 480954 554614 481574 576000
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 466308 481574 482058
rect 487794 561454 488414 576000
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 466308 488414 488898
rect 488582 486437 488642 627811
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 491514 565174 492134 576000
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 488579 486436 488645 486437
rect 488579 486372 488580 486436
rect 488644 486372 488645 486436
rect 488579 486371 488645 486372
rect 491514 466308 492134 492618
rect 495234 568894 495854 576000
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 466308 495854 496338
rect 498954 572614 499574 576000
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498515 466580 498581 466581
rect 498515 466516 498516 466580
rect 498580 466516 498581 466580
rect 498515 466515 498581 466516
rect 498518 464810 498578 466515
rect 498954 466308 499574 500058
rect 505794 543454 506414 576000
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 506614 472701 506674 627811
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 509514 547174 510134 576000
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 506611 472700 506677 472701
rect 506611 472636 506612 472700
rect 506676 472636 506677 472700
rect 506611 472635 506677 472636
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 499803 466580 499869 466581
rect 499803 466516 499804 466580
rect 499868 466516 499869 466580
rect 499803 466515 499869 466516
rect 499806 464810 499866 466515
rect 505794 466308 506414 470898
rect 509514 466308 510134 474618
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 510843 466580 510909 466581
rect 510843 466516 510844 466580
rect 510908 466516 510909 466580
rect 510843 466515 510909 466516
rect 510846 464810 510906 466515
rect 513234 466308 513854 478338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 466308 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 498464 464750 498578 464810
rect 499688 464750 499866 464810
rect 510840 464750 510906 464810
rect 498464 464202 498524 464750
rect 499688 464202 499748 464750
rect 510840 464202 510900 464750
rect 380272 453454 380620 453486
rect 380272 453218 380328 453454
rect 380564 453218 380620 453454
rect 380272 453134 380620 453218
rect 380272 452898 380328 453134
rect 380564 452898 380620 453134
rect 380272 452866 380620 452898
rect 516000 453454 516348 453486
rect 516000 453218 516056 453454
rect 516292 453218 516348 453454
rect 516000 453134 516348 453218
rect 516000 452898 516056 453134
rect 516292 452898 516348 453134
rect 516000 452866 516348 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 380952 435454 381300 435486
rect 380952 435218 381008 435454
rect 381244 435218 381300 435454
rect 380952 435134 381300 435218
rect 380952 434898 381008 435134
rect 381244 434898 381300 435134
rect 380952 434866 381300 434898
rect 515320 435454 515668 435486
rect 515320 435218 515376 435454
rect 515612 435218 515668 435454
rect 515320 435134 515668 435218
rect 515320 434898 515376 435134
rect 515612 434898 515668 435134
rect 515320 434866 515668 434898
rect 380272 417454 380620 417486
rect 380272 417218 380328 417454
rect 380564 417218 380620 417454
rect 380272 417134 380620 417218
rect 380272 416898 380328 417134
rect 380564 416898 380620 417134
rect 380272 416866 380620 416898
rect 516000 417454 516348 417486
rect 516000 417218 516056 417454
rect 516292 417218 516348 417454
rect 516000 417134 516348 417218
rect 516000 416898 516056 417134
rect 516292 416898 516348 417134
rect 516000 416866 516348 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 380952 399454 381300 399486
rect 380952 399218 381008 399454
rect 381244 399218 381300 399454
rect 380952 399134 381300 399218
rect 380952 398898 381008 399134
rect 381244 398898 381300 399134
rect 380952 398866 381300 398898
rect 515320 399454 515668 399486
rect 515320 399218 515376 399454
rect 515612 399218 515668 399454
rect 515320 399134 515668 399218
rect 515320 398898 515376 399134
rect 515612 398898 515668 399134
rect 515320 398866 515668 398898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 396056 380490 396116 381106
rect 397144 380490 397204 381106
rect 396030 380430 396116 380490
rect 397134 380430 397204 380490
rect 398232 380490 398292 381106
rect 399592 380490 399652 381106
rect 400544 380490 400604 381106
rect 398232 380430 398298 380490
rect 396030 379405 396090 380430
rect 397134 379405 397194 380430
rect 396027 379404 396093 379405
rect 396027 379340 396028 379404
rect 396092 379340 396093 379404
rect 396027 379339 396093 379340
rect 397131 379404 397197 379405
rect 397131 379340 397132 379404
rect 397196 379340 397197 379404
rect 397131 379339 397197 379340
rect 398238 379269 398298 380430
rect 399526 380430 399652 380490
rect 400446 380430 400604 380490
rect 401768 380490 401828 381106
rect 403128 380490 403188 381106
rect 404216 380490 404276 381106
rect 405440 380490 405500 381106
rect 406528 380490 406588 381106
rect 401768 380430 402346 380490
rect 398235 379268 398301 379269
rect 398235 379204 398236 379268
rect 398300 379204 398301 379268
rect 398235 379203 398301 379204
rect 399526 379133 399586 380430
rect 399523 379132 399589 379133
rect 399523 379068 399524 379132
rect 399588 379068 399589 379132
rect 399523 379067 399589 379068
rect 379794 364394 380414 379000
rect 379794 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 380414 364394
rect 379794 364074 380414 364158
rect 379794 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 380414 364074
rect 379794 359308 380414 363838
rect 383514 368114 384134 379000
rect 383514 367878 383546 368114
rect 383782 367878 383866 368114
rect 384102 367878 384134 368114
rect 383514 367794 384134 367878
rect 383514 367558 383546 367794
rect 383782 367558 383866 367794
rect 384102 367558 384134 367794
rect 383514 359308 384134 367558
rect 387234 369954 387854 379000
rect 387234 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 387854 369954
rect 387234 369634 387854 369718
rect 387234 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 387854 369634
rect 387234 359308 387854 369398
rect 390954 373674 391574 379000
rect 390954 373438 390986 373674
rect 391222 373438 391306 373674
rect 391542 373438 391574 373674
rect 390954 373354 391574 373438
rect 390954 373118 390986 373354
rect 391222 373118 391306 373354
rect 391542 373118 391574 373354
rect 390954 359308 391574 373118
rect 397794 363454 398414 379000
rect 400446 378725 400506 380430
rect 400443 378724 400509 378725
rect 400443 378660 400444 378724
rect 400508 378660 400509 378724
rect 400443 378659 400509 378660
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 359308 398414 362898
rect 401514 367174 402134 379000
rect 402286 378861 402346 380430
rect 403022 380430 403188 380490
rect 404126 380430 404276 380490
rect 405414 380430 405500 380490
rect 406518 380430 406588 380490
rect 407616 380490 407676 381106
rect 408296 380490 408356 381106
rect 408704 380629 408764 381106
rect 408701 380628 408767 380629
rect 408701 380564 408702 380628
rect 408766 380564 408767 380628
rect 408701 380563 408767 380564
rect 410064 380490 410124 381106
rect 407616 380430 407682 380490
rect 408296 380430 408418 380490
rect 403022 379269 403082 380430
rect 404126 379405 404186 380430
rect 404123 379404 404189 379405
rect 404123 379340 404124 379404
rect 404188 379340 404189 379404
rect 404123 379339 404189 379340
rect 405414 379269 405474 380430
rect 406518 379405 406578 380430
rect 407622 379405 407682 380430
rect 408358 379405 408418 380430
rect 410014 380430 410124 380490
rect 410744 380490 410804 381106
rect 411288 380490 411348 381106
rect 412376 380490 412436 381106
rect 413464 380629 413524 381106
rect 413461 380628 413527 380629
rect 413461 380564 413462 380628
rect 413526 380564 413527 380628
rect 413461 380563 413527 380564
rect 413600 380490 413660 381106
rect 410744 380430 410810 380490
rect 411288 380430 411362 380490
rect 412376 380430 412466 380490
rect 406515 379404 406581 379405
rect 406515 379340 406516 379404
rect 406580 379340 406581 379404
rect 406515 379339 406581 379340
rect 407619 379404 407685 379405
rect 407619 379340 407620 379404
rect 407684 379340 407685 379404
rect 407619 379339 407685 379340
rect 408355 379404 408421 379405
rect 408355 379340 408356 379404
rect 408420 379340 408421 379404
rect 408355 379339 408421 379340
rect 403019 379268 403085 379269
rect 403019 379204 403020 379268
rect 403084 379204 403085 379268
rect 403019 379203 403085 379204
rect 405411 379268 405477 379269
rect 405411 379204 405412 379268
rect 405476 379204 405477 379268
rect 405411 379203 405477 379204
rect 402283 378860 402349 378861
rect 402283 378796 402284 378860
rect 402348 378796 402349 378860
rect 402283 378795 402349 378796
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 359308 402134 366618
rect 405234 370894 405854 379000
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 359308 405854 370338
rect 408954 374614 409574 379000
rect 410014 378181 410074 380430
rect 410750 379269 410810 380430
rect 411302 379405 411362 380430
rect 412406 379405 412466 380430
rect 413510 380430 413660 380490
rect 414552 380490 414612 381106
rect 415912 380490 415972 381106
rect 414552 380430 414674 380490
rect 413510 379405 413570 380430
rect 414614 379405 414674 380430
rect 415902 380430 415972 380490
rect 416048 380490 416108 381106
rect 417000 380490 417060 381106
rect 418088 380490 418148 381106
rect 418496 380490 418556 381106
rect 419448 380629 419508 381106
rect 419445 380628 419511 380629
rect 419445 380564 419446 380628
rect 419510 380564 419511 380628
rect 419445 380563 419511 380564
rect 416048 380430 416146 380490
rect 417000 380430 417066 380490
rect 418088 380430 418170 380490
rect 411299 379404 411365 379405
rect 411299 379340 411300 379404
rect 411364 379340 411365 379404
rect 411299 379339 411365 379340
rect 412403 379404 412469 379405
rect 412403 379340 412404 379404
rect 412468 379340 412469 379404
rect 412403 379339 412469 379340
rect 413507 379404 413573 379405
rect 413507 379340 413508 379404
rect 413572 379340 413573 379404
rect 413507 379339 413573 379340
rect 414611 379404 414677 379405
rect 414611 379340 414612 379404
rect 414676 379340 414677 379404
rect 414611 379339 414677 379340
rect 415902 379269 415962 380430
rect 416086 379269 416146 380430
rect 410747 379268 410813 379269
rect 410747 379204 410748 379268
rect 410812 379204 410813 379268
rect 410747 379203 410813 379204
rect 415899 379268 415965 379269
rect 415899 379204 415900 379268
rect 415964 379204 415965 379268
rect 415899 379203 415965 379204
rect 416083 379268 416149 379269
rect 416083 379204 416084 379268
rect 416148 379204 416149 379268
rect 416083 379203 416149 379204
rect 410011 378180 410077 378181
rect 410011 378116 410012 378180
rect 410076 378116 410077 378180
rect 410011 378115 410077 378116
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 359308 409574 374058
rect 415794 364394 416414 379000
rect 417006 378589 417066 380430
rect 417003 378588 417069 378589
rect 417003 378524 417004 378588
rect 417068 378524 417069 378588
rect 417003 378523 417069 378524
rect 418110 378181 418170 380430
rect 418478 380430 418556 380490
rect 420672 380490 420732 381106
rect 421080 380765 421140 381106
rect 421077 380764 421143 380765
rect 421077 380700 421078 380764
rect 421142 380700 421143 380764
rect 421077 380699 421143 380700
rect 421760 380490 421820 381106
rect 422848 380765 422908 381106
rect 422845 380764 422911 380765
rect 422845 380700 422846 380764
rect 422910 380700 422911 380764
rect 422845 380699 422911 380700
rect 423528 380490 423588 381106
rect 420672 380430 420746 380490
rect 421760 380430 421850 380490
rect 418478 378725 418538 380430
rect 418475 378724 418541 378725
rect 418475 378660 418476 378724
rect 418540 378660 418541 378724
rect 418475 378659 418541 378660
rect 418107 378180 418173 378181
rect 418107 378116 418108 378180
rect 418172 378116 418173 378180
rect 418107 378115 418173 378116
rect 415794 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 416414 364394
rect 415794 364074 416414 364158
rect 415794 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 416414 364074
rect 415794 359308 416414 363838
rect 419514 368114 420134 379000
rect 420686 378181 420746 380430
rect 421790 378181 421850 380430
rect 423446 380430 423588 380490
rect 423936 380490 423996 381106
rect 425296 380490 425356 381106
rect 423936 380430 424058 380490
rect 423446 379405 423506 380430
rect 423443 379404 423509 379405
rect 423443 379340 423444 379404
rect 423508 379340 423509 379404
rect 423443 379339 423509 379340
rect 420683 378180 420749 378181
rect 420683 378116 420684 378180
rect 420748 378116 420749 378180
rect 420683 378115 420749 378116
rect 421787 378180 421853 378181
rect 421787 378116 421788 378180
rect 421852 378116 421853 378180
rect 421787 378115 421853 378116
rect 419514 367878 419546 368114
rect 419782 367878 419866 368114
rect 420102 367878 420134 368114
rect 419514 367794 420134 367878
rect 419514 367558 419546 367794
rect 419782 367558 419866 367794
rect 420102 367558 420134 367794
rect 419514 359308 420134 367558
rect 423234 369954 423854 379000
rect 423998 378181 424058 380430
rect 425286 380430 425356 380490
rect 425976 380490 426036 381106
rect 426384 380490 426444 381106
rect 427608 380490 427668 381106
rect 428288 380490 428348 381106
rect 428696 380490 428756 381106
rect 429784 380490 429844 381106
rect 431008 380765 431068 381106
rect 431005 380764 431071 380765
rect 431005 380700 431006 380764
rect 431070 380700 431071 380764
rect 431005 380699 431071 380700
rect 425976 380430 426082 380490
rect 426384 380430 426450 380490
rect 425286 378181 425346 380430
rect 426022 378725 426082 380430
rect 426390 379405 426450 380430
rect 427494 380430 427668 380490
rect 428230 380430 428348 380490
rect 428598 380430 428756 380490
rect 429702 380430 429844 380490
rect 431144 380490 431204 381106
rect 432232 380490 432292 381106
rect 433320 380490 433380 381106
rect 433592 380765 433652 381106
rect 433589 380764 433655 380765
rect 433589 380700 433590 380764
rect 433654 380700 433655 380764
rect 433589 380699 433655 380700
rect 434408 380629 434468 381106
rect 434405 380628 434471 380629
rect 434405 380564 434406 380628
rect 434470 380564 434471 380628
rect 434405 380563 434471 380564
rect 435768 380490 435828 381106
rect 436040 380765 436100 381106
rect 436037 380764 436103 380765
rect 436037 380700 436038 380764
rect 436102 380700 436103 380764
rect 436037 380699 436103 380700
rect 436992 380490 437052 381106
rect 438080 380490 438140 381106
rect 438488 380765 438548 381106
rect 438485 380764 438551 380765
rect 438485 380700 438486 380764
rect 438550 380700 438551 380764
rect 438485 380699 438551 380700
rect 439168 380490 439228 381106
rect 440936 380765 440996 381106
rect 443520 380765 443580 381106
rect 440933 380764 440999 380765
rect 440933 380700 440934 380764
rect 440998 380700 440999 380764
rect 440933 380699 440999 380700
rect 443517 380764 443583 380765
rect 443517 380700 443518 380764
rect 443582 380700 443583 380764
rect 443517 380699 443583 380700
rect 445968 380629 446028 381106
rect 445965 380628 446031 380629
rect 445965 380564 445966 380628
rect 446030 380564 446031 380628
rect 445965 380563 446031 380564
rect 431144 380430 431234 380490
rect 432232 380430 432338 380490
rect 433320 380430 433442 380490
rect 435768 380430 435834 380490
rect 427494 379405 427554 380430
rect 426387 379404 426453 379405
rect 426387 379340 426388 379404
rect 426452 379340 426453 379404
rect 426387 379339 426453 379340
rect 427491 379404 427557 379405
rect 427491 379340 427492 379404
rect 427556 379340 427557 379404
rect 427491 379339 427557 379340
rect 426019 378724 426085 378725
rect 426019 378660 426020 378724
rect 426084 378660 426085 378724
rect 426019 378659 426085 378660
rect 423995 378180 424061 378181
rect 423995 378116 423996 378180
rect 424060 378116 424061 378180
rect 423995 378115 424061 378116
rect 425283 378180 425349 378181
rect 425283 378116 425284 378180
rect 425348 378116 425349 378180
rect 425283 378115 425349 378116
rect 423234 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 423854 369954
rect 423234 369634 423854 369718
rect 423234 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 423854 369634
rect 423234 359308 423854 369398
rect 426954 373674 427574 379000
rect 428230 378725 428290 380430
rect 428227 378724 428293 378725
rect 428227 378660 428228 378724
rect 428292 378660 428293 378724
rect 428227 378659 428293 378660
rect 428598 378181 428658 380430
rect 429702 378181 429762 380430
rect 431174 378317 431234 380430
rect 431171 378316 431237 378317
rect 431171 378252 431172 378316
rect 431236 378252 431237 378316
rect 431171 378251 431237 378252
rect 432278 378181 432338 380430
rect 433382 379133 433442 380430
rect 435774 379405 435834 380430
rect 436878 380430 437052 380490
rect 437982 380430 438140 380490
rect 439086 380430 439228 380490
rect 448280 380490 448340 381106
rect 451000 380490 451060 381106
rect 453448 380490 453508 381106
rect 455896 380490 455956 381106
rect 458480 380490 458540 381106
rect 448280 380430 448346 380490
rect 451000 380430 451106 380490
rect 435771 379404 435837 379405
rect 435771 379340 435772 379404
rect 435836 379340 435837 379404
rect 435771 379339 435837 379340
rect 433379 379132 433445 379133
rect 433379 379068 433380 379132
rect 433444 379068 433445 379132
rect 433379 379067 433445 379068
rect 428595 378180 428661 378181
rect 428595 378116 428596 378180
rect 428660 378116 428661 378180
rect 428595 378115 428661 378116
rect 429699 378180 429765 378181
rect 429699 378116 429700 378180
rect 429764 378116 429765 378180
rect 429699 378115 429765 378116
rect 432275 378180 432341 378181
rect 432275 378116 432276 378180
rect 432340 378116 432341 378180
rect 432275 378115 432341 378116
rect 426954 373438 426986 373674
rect 427222 373438 427306 373674
rect 427542 373438 427574 373674
rect 426954 373354 427574 373438
rect 426954 373118 426986 373354
rect 427222 373118 427306 373354
rect 427542 373118 427574 373354
rect 426954 359308 427574 373118
rect 433794 363454 434414 379000
rect 436878 378589 436938 380430
rect 437982 379269 438042 380430
rect 439086 379405 439146 380430
rect 448286 379405 448346 380430
rect 451046 379405 451106 380430
rect 453438 380430 453508 380490
rect 455830 380430 455956 380490
rect 458406 380430 458540 380490
rect 460928 380490 460988 381106
rect 463512 380490 463572 381106
rect 465960 380490 466020 381106
rect 468544 380490 468604 381106
rect 470992 380490 471052 381106
rect 460928 380430 461042 380490
rect 463512 380430 463618 380490
rect 453438 379405 453498 380430
rect 455830 379405 455890 380430
rect 458406 379405 458466 380430
rect 460982 379405 461042 380430
rect 463558 379405 463618 380430
rect 465950 380430 466020 380490
rect 468526 380430 468604 380490
rect 470918 380430 471052 380490
rect 473440 380490 473500 381106
rect 475888 380490 475948 381106
rect 478472 380490 478532 381106
rect 480920 380490 480980 381106
rect 473440 380430 473554 380490
rect 439083 379404 439149 379405
rect 439083 379340 439084 379404
rect 439148 379340 439149 379404
rect 439083 379339 439149 379340
rect 448283 379404 448349 379405
rect 448283 379340 448284 379404
rect 448348 379340 448349 379404
rect 448283 379339 448349 379340
rect 451043 379404 451109 379405
rect 451043 379340 451044 379404
rect 451108 379340 451109 379404
rect 451043 379339 451109 379340
rect 453435 379404 453501 379405
rect 453435 379340 453436 379404
rect 453500 379340 453501 379404
rect 453435 379339 453501 379340
rect 455827 379404 455893 379405
rect 455827 379340 455828 379404
rect 455892 379340 455893 379404
rect 455827 379339 455893 379340
rect 458403 379404 458469 379405
rect 458403 379340 458404 379404
rect 458468 379340 458469 379404
rect 458403 379339 458469 379340
rect 460979 379404 461045 379405
rect 460979 379340 460980 379404
rect 461044 379340 461045 379404
rect 460979 379339 461045 379340
rect 463555 379404 463621 379405
rect 463555 379340 463556 379404
rect 463620 379340 463621 379404
rect 463555 379339 463621 379340
rect 437979 379268 438045 379269
rect 437979 379204 437980 379268
rect 438044 379204 438045 379268
rect 437979 379203 438045 379204
rect 465950 379133 466010 380430
rect 465947 379132 466013 379133
rect 465947 379068 465948 379132
rect 466012 379068 466013 379132
rect 465947 379067 466013 379068
rect 436875 378588 436941 378589
rect 436875 378524 436876 378588
rect 436940 378524 436941 378588
rect 436875 378523 436941 378524
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 359308 434414 362898
rect 437514 367174 438134 379000
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 359308 438134 366618
rect 441234 370894 441854 379000
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 359308 441854 370338
rect 444954 374614 445574 379000
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 359308 445574 374058
rect 451794 364394 452414 379000
rect 451794 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 452414 364394
rect 451794 364074 452414 364158
rect 451794 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 452414 364074
rect 451794 359308 452414 363838
rect 455514 368114 456134 379000
rect 455514 367878 455546 368114
rect 455782 367878 455866 368114
rect 456102 367878 456134 368114
rect 455514 367794 456134 367878
rect 455514 367558 455546 367794
rect 455782 367558 455866 367794
rect 456102 367558 456134 367794
rect 455514 359308 456134 367558
rect 459234 369954 459854 379000
rect 459234 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 459854 369954
rect 459234 369634 459854 369718
rect 459234 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 459854 369634
rect 459234 359308 459854 369398
rect 462954 373674 463574 379000
rect 468526 378861 468586 380430
rect 468523 378860 468589 378861
rect 468523 378796 468524 378860
rect 468588 378796 468589 378860
rect 468523 378795 468589 378796
rect 462954 373438 462986 373674
rect 463222 373438 463306 373674
rect 463542 373438 463574 373674
rect 462954 373354 463574 373438
rect 462954 373118 462986 373354
rect 463222 373118 463306 373354
rect 463542 373118 463574 373354
rect 462954 359308 463574 373118
rect 469794 363454 470414 379000
rect 470918 378861 470978 380430
rect 473494 379269 473554 380430
rect 475886 380430 475948 380490
rect 478462 380430 478532 380490
rect 480854 380430 480980 380490
rect 483368 380490 483428 381106
rect 485952 380901 486012 381106
rect 485949 380900 486015 380901
rect 485949 380836 485950 380900
rect 486014 380836 486015 380900
rect 485949 380835 486015 380836
rect 503224 380490 503284 381106
rect 483368 380430 483490 380490
rect 475886 379405 475946 380430
rect 475883 379404 475949 379405
rect 475883 379340 475884 379404
rect 475948 379340 475949 379404
rect 475883 379339 475949 379340
rect 473491 379268 473557 379269
rect 473491 379204 473492 379268
rect 473556 379204 473557 379268
rect 473491 379203 473557 379204
rect 470915 378860 470981 378861
rect 470915 378796 470916 378860
rect 470980 378796 470981 378860
rect 470915 378795 470981 378796
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 359308 470414 362898
rect 473514 367174 474134 379000
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 359308 474134 366618
rect 477234 370894 477854 379000
rect 478462 378997 478522 380430
rect 480854 379269 480914 380430
rect 480851 379268 480917 379269
rect 480851 379204 480852 379268
rect 480916 379204 480917 379268
rect 480851 379203 480917 379204
rect 478459 378996 478525 378997
rect 478459 378932 478460 378996
rect 478524 378932 478525 378996
rect 478459 378931 478525 378932
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 359308 477854 370338
rect 480954 374614 481574 379000
rect 483430 378997 483490 380430
rect 503118 380430 503284 380490
rect 503360 380490 503420 381106
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 503360 380430 503546 380490
rect 503118 379269 503178 380430
rect 503486 379269 503546 380430
rect 503115 379268 503181 379269
rect 503115 379204 503116 379268
rect 503180 379204 503181 379268
rect 503115 379203 503181 379204
rect 503483 379268 503549 379269
rect 503483 379204 503484 379268
rect 503548 379204 503549 379268
rect 503483 379203 503549 379204
rect 483427 378996 483493 378997
rect 483427 378932 483428 378996
rect 483492 378932 483493 378996
rect 483427 378931 483493 378932
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 359308 481574 374058
rect 487794 364394 488414 379000
rect 487794 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 487794 364074 488414 364158
rect 487794 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 487794 359308 488414 363838
rect 491514 368114 492134 379000
rect 491514 367878 491546 368114
rect 491782 367878 491866 368114
rect 492102 367878 492134 368114
rect 491514 367794 492134 367878
rect 491514 367558 491546 367794
rect 491782 367558 491866 367794
rect 492102 367558 492134 367794
rect 491514 359308 492134 367558
rect 495234 369954 495854 379000
rect 495234 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 495234 369634 495854 369718
rect 495234 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 495234 359308 495854 369398
rect 498954 373674 499574 379000
rect 498954 373438 498986 373674
rect 499222 373438 499306 373674
rect 499542 373438 499574 373674
rect 498954 373354 499574 373438
rect 498954 373118 498986 373354
rect 499222 373118 499306 373354
rect 499542 373118 499574 373354
rect 498954 359308 499574 373118
rect 505794 363454 506414 379000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 359308 506414 362898
rect 509514 367174 510134 379000
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 359308 510134 366618
rect 513234 370894 513854 379000
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 359308 513854 370338
rect 516954 374614 517574 379000
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 359308 517574 374058
rect 498515 358868 498581 358869
rect 498515 358804 498516 358868
rect 498580 358804 498581 358868
rect 498515 358803 498581 358804
rect 499803 358868 499869 358869
rect 499803 358804 499804 358868
rect 499868 358804 499869 358868
rect 499803 358803 499869 358804
rect 510843 358868 510909 358869
rect 510843 358804 510844 358868
rect 510908 358804 510909 358868
rect 510843 358803 510909 358804
rect 498518 358050 498578 358803
rect 499806 358050 499866 358803
rect 510846 358050 510906 358803
rect 498464 357990 498578 358050
rect 499688 357990 499866 358050
rect 510840 357990 510906 358050
rect 498464 357202 498524 357990
rect 499688 357202 499748 357990
rect 510840 357202 510900 357990
rect 380272 345454 380620 345486
rect 380272 345218 380328 345454
rect 380564 345218 380620 345454
rect 380272 345134 380620 345218
rect 380272 344898 380328 345134
rect 380564 344898 380620 345134
rect 380272 344866 380620 344898
rect 516000 345454 516348 345486
rect 516000 345218 516056 345454
rect 516292 345218 516348 345454
rect 516000 345134 516348 345218
rect 516000 344898 516056 345134
rect 516292 344898 516348 345134
rect 516000 344866 516348 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 380952 327454 381300 327486
rect 380952 327218 381008 327454
rect 381244 327218 381300 327454
rect 380952 327134 381300 327218
rect 380952 326898 381008 327134
rect 381244 326898 381300 327134
rect 380952 326866 381300 326898
rect 515320 327454 515668 327486
rect 515320 327218 515376 327454
rect 515612 327218 515668 327454
rect 515320 327134 515668 327218
rect 515320 326898 515376 327134
rect 515612 326898 515668 327134
rect 515320 326866 515668 326898
rect 380272 309454 380620 309486
rect 380272 309218 380328 309454
rect 380564 309218 380620 309454
rect 380272 309134 380620 309218
rect 380272 308898 380328 309134
rect 380564 308898 380620 309134
rect 380272 308866 380620 308898
rect 516000 309454 516348 309486
rect 516000 309218 516056 309454
rect 516292 309218 516348 309454
rect 516000 309134 516348 309218
rect 516000 308898 516056 309134
rect 516292 308898 516348 309134
rect 516000 308866 516348 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 380952 291454 381300 291486
rect 380952 291218 381008 291454
rect 381244 291218 381300 291454
rect 380952 291134 381300 291218
rect 380952 290898 381008 291134
rect 381244 290898 381300 291134
rect 380952 290866 381300 290898
rect 515320 291454 515668 291486
rect 515320 291218 515376 291454
rect 515612 291218 515668 291454
rect 515320 291134 515668 291218
rect 515320 290898 515376 291134
rect 515612 290898 515668 291134
rect 515320 290866 515668 290898
rect 396056 273730 396116 274040
rect 397144 273730 397204 274040
rect 398232 273730 398292 274040
rect 399592 273730 399652 274040
rect 400544 273730 400604 274040
rect 401768 273730 401828 274040
rect 403128 273730 403188 274040
rect 404216 273730 404276 274040
rect 405440 273730 405500 274040
rect 406528 273730 406588 274040
rect 396030 273670 396116 273730
rect 397134 273670 397204 273730
rect 397502 273670 398292 273730
rect 399526 273670 399652 273730
rect 400446 273670 400604 273730
rect 401734 273670 401828 273730
rect 403022 273670 403188 273730
rect 404126 273670 404276 273730
rect 405046 273670 405500 273730
rect 406518 273670 406588 273730
rect 407616 273730 407676 274040
rect 408296 273730 408356 274040
rect 407616 273670 407682 273730
rect 379794 256394 380414 272000
rect 379794 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 380414 256394
rect 379794 256074 380414 256158
rect 379794 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 380414 256074
rect 379794 252308 380414 255838
rect 383514 260114 384134 272000
rect 383514 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 384134 260114
rect 383514 259794 384134 259878
rect 383514 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 384134 259794
rect 383514 252308 384134 259558
rect 387234 261954 387854 272000
rect 387234 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 387854 261954
rect 387234 261634 387854 261718
rect 387234 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 387854 261634
rect 387234 252308 387854 261398
rect 390954 265674 391574 272000
rect 396030 271285 396090 273670
rect 396027 271284 396093 271285
rect 396027 271220 396028 271284
rect 396092 271220 396093 271284
rect 396027 271219 396093 271220
rect 397134 271149 397194 273670
rect 397131 271148 397197 271149
rect 397131 271084 397132 271148
rect 397196 271084 397197 271148
rect 397131 271083 397197 271084
rect 397502 270605 397562 273670
rect 397499 270604 397565 270605
rect 397499 270540 397500 270604
rect 397564 270540 397565 270604
rect 397499 270539 397565 270540
rect 390954 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 391574 265674
rect 390954 265354 391574 265438
rect 390954 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 391574 265354
rect 390954 252308 391574 265118
rect 397794 255454 398414 272000
rect 399526 270605 399586 273670
rect 400446 270605 400506 273670
rect 401734 272237 401794 273670
rect 401731 272236 401797 272237
rect 401731 272172 401732 272236
rect 401796 272172 401797 272236
rect 401731 272171 401797 272172
rect 399523 270604 399589 270605
rect 399523 270540 399524 270604
rect 399588 270540 399589 270604
rect 399523 270539 399589 270540
rect 400443 270604 400509 270605
rect 400443 270540 400444 270604
rect 400508 270540 400509 270604
rect 400443 270539 400509 270540
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 252308 398414 254898
rect 401514 259174 402134 272000
rect 403022 270605 403082 273670
rect 404126 270605 404186 273670
rect 405046 270605 405106 273670
rect 403019 270604 403085 270605
rect 403019 270540 403020 270604
rect 403084 270540 403085 270604
rect 403019 270539 403085 270540
rect 404123 270604 404189 270605
rect 404123 270540 404124 270604
rect 404188 270540 404189 270604
rect 404123 270539 404189 270540
rect 405043 270604 405109 270605
rect 405043 270540 405044 270604
rect 405108 270540 405109 270604
rect 405043 270539 405109 270540
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 252308 402134 258618
rect 405234 262894 405854 272000
rect 406518 270877 406578 273670
rect 406515 270876 406581 270877
rect 406515 270812 406516 270876
rect 406580 270812 406581 270876
rect 406515 270811 406581 270812
rect 407622 270605 407682 273670
rect 408174 273670 408356 273730
rect 408704 273730 408764 274040
rect 410064 273730 410124 274040
rect 408704 273670 408786 273730
rect 408174 271421 408234 273670
rect 408171 271420 408237 271421
rect 408171 271356 408172 271420
rect 408236 271356 408237 271420
rect 408171 271355 408237 271356
rect 408726 270605 408786 273670
rect 410014 273670 410124 273730
rect 410744 273730 410804 274040
rect 411288 273730 411348 274040
rect 412376 273730 412436 274040
rect 413464 273730 413524 274040
rect 410744 273670 410810 273730
rect 411288 273670 411362 273730
rect 412376 273670 412466 273730
rect 407619 270604 407685 270605
rect 407619 270540 407620 270604
rect 407684 270540 407685 270604
rect 407619 270539 407685 270540
rect 408723 270604 408789 270605
rect 408723 270540 408724 270604
rect 408788 270540 408789 270604
rect 408723 270539 408789 270540
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 252308 405854 262338
rect 408954 266614 409574 272000
rect 410014 270605 410074 273670
rect 410750 271149 410810 273670
rect 410747 271148 410813 271149
rect 410747 271084 410748 271148
rect 410812 271084 410813 271148
rect 410747 271083 410813 271084
rect 411302 270741 411362 273670
rect 411299 270740 411365 270741
rect 411299 270676 411300 270740
rect 411364 270676 411365 270740
rect 411299 270675 411365 270676
rect 412406 270605 412466 273670
rect 413326 273670 413524 273730
rect 413600 273730 413660 274040
rect 414552 273730 414612 274040
rect 415912 273730 415972 274040
rect 413600 273670 413754 273730
rect 413326 270605 413386 273670
rect 413694 271149 413754 273670
rect 414430 273670 414612 273730
rect 415902 273670 415972 273730
rect 416048 273730 416108 274040
rect 417000 273730 417060 274040
rect 418088 273730 418148 274040
rect 418496 273730 418556 274040
rect 419448 273730 419508 274040
rect 416048 273670 416146 273730
rect 417000 273670 417066 273730
rect 418088 273670 418170 273730
rect 413691 271148 413757 271149
rect 413691 271084 413692 271148
rect 413756 271084 413757 271148
rect 413691 271083 413757 271084
rect 414430 270605 414490 273670
rect 415902 272237 415962 273670
rect 416086 272237 416146 273670
rect 415899 272236 415965 272237
rect 415899 272172 415900 272236
rect 415964 272172 415965 272236
rect 415899 272171 415965 272172
rect 416083 272236 416149 272237
rect 416083 272172 416084 272236
rect 416148 272172 416149 272236
rect 416083 272171 416149 272172
rect 410011 270604 410077 270605
rect 410011 270540 410012 270604
rect 410076 270540 410077 270604
rect 410011 270539 410077 270540
rect 412403 270604 412469 270605
rect 412403 270540 412404 270604
rect 412468 270540 412469 270604
rect 412403 270539 412469 270540
rect 413323 270604 413389 270605
rect 413323 270540 413324 270604
rect 413388 270540 413389 270604
rect 413323 270539 413389 270540
rect 414427 270604 414493 270605
rect 414427 270540 414428 270604
rect 414492 270540 414493 270604
rect 414427 270539 414493 270540
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 252308 409574 266058
rect 415794 256394 416414 272000
rect 417006 270605 417066 273670
rect 418110 270605 418170 273670
rect 418478 273670 418556 273730
rect 419214 273670 419508 273730
rect 420672 273730 420732 274040
rect 420672 273670 420746 273730
rect 418478 271149 418538 273670
rect 418475 271148 418541 271149
rect 418475 271084 418476 271148
rect 418540 271084 418541 271148
rect 418475 271083 418541 271084
rect 417003 270604 417069 270605
rect 417003 270540 417004 270604
rect 417068 270540 417069 270604
rect 417003 270539 417069 270540
rect 418107 270604 418173 270605
rect 418107 270540 418108 270604
rect 418172 270540 418173 270604
rect 418107 270539 418173 270540
rect 419214 270469 419274 273670
rect 419211 270468 419277 270469
rect 419211 270404 419212 270468
rect 419276 270404 419277 270468
rect 419211 270403 419277 270404
rect 415794 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 416414 256394
rect 415794 256074 416414 256158
rect 415794 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 416414 256074
rect 415794 252308 416414 255838
rect 419514 260114 420134 272000
rect 420686 270605 420746 273670
rect 421080 273597 421140 274040
rect 421760 273730 421820 274040
rect 421760 273670 421850 273730
rect 421077 273596 421143 273597
rect 421077 273532 421078 273596
rect 421142 273532 421143 273596
rect 421077 273531 421143 273532
rect 421790 270605 421850 273670
rect 422848 273597 422908 274040
rect 423528 273730 423588 274040
rect 423936 273730 423996 274040
rect 425296 273730 425356 274040
rect 423446 273670 423588 273730
rect 423814 273670 423996 273730
rect 425286 273670 425356 273730
rect 425976 273730 426036 274040
rect 426384 273730 426444 274040
rect 425976 273670 426082 273730
rect 426384 273670 426450 273730
rect 422845 273596 422911 273597
rect 422845 273532 422846 273596
rect 422910 273532 422911 273596
rect 422845 273531 422911 273532
rect 423446 273053 423506 273670
rect 423443 273052 423509 273053
rect 423443 272988 423444 273052
rect 423508 272988 423509 273052
rect 423443 272987 423509 272988
rect 423814 272917 423874 273670
rect 425286 273053 425346 273670
rect 426022 273053 426082 273670
rect 425283 273052 425349 273053
rect 425283 272988 425284 273052
rect 425348 272988 425349 273052
rect 425283 272987 425349 272988
rect 426019 273052 426085 273053
rect 426019 272988 426020 273052
rect 426084 272988 426085 273052
rect 426019 272987 426085 272988
rect 423811 272916 423877 272917
rect 423811 272852 423812 272916
rect 423876 272852 423877 272916
rect 423811 272851 423877 272852
rect 420683 270604 420749 270605
rect 420683 270540 420684 270604
rect 420748 270540 420749 270604
rect 420683 270539 420749 270540
rect 421787 270604 421853 270605
rect 421787 270540 421788 270604
rect 421852 270540 421853 270604
rect 421787 270539 421853 270540
rect 419514 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 420134 260114
rect 419514 259794 420134 259878
rect 419514 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 420134 259794
rect 419514 252308 420134 259558
rect 423234 261954 423854 272000
rect 426390 269789 426450 273670
rect 427608 273597 427668 274040
rect 428288 273730 428348 274040
rect 428696 273730 428756 274040
rect 429784 273730 429844 274040
rect 431008 273730 431068 274040
rect 428230 273670 428348 273730
rect 428598 273670 428756 273730
rect 429702 273670 429844 273730
rect 430990 273670 431068 273730
rect 431144 273730 431204 274040
rect 432232 273730 432292 274040
rect 433320 273730 433380 274040
rect 433592 273730 433652 274040
rect 431144 273670 431234 273730
rect 432232 273670 432338 273730
rect 433320 273670 433442 273730
rect 427605 273596 427671 273597
rect 427605 273532 427606 273596
rect 427670 273532 427671 273596
rect 427605 273531 427671 273532
rect 428230 273053 428290 273670
rect 428227 273052 428293 273053
rect 428227 272988 428228 273052
rect 428292 272988 428293 273052
rect 428227 272987 428293 272988
rect 426387 269788 426453 269789
rect 426387 269724 426388 269788
rect 426452 269724 426453 269788
rect 426387 269723 426453 269724
rect 423234 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 423854 261954
rect 423234 261634 423854 261718
rect 423234 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 423854 261634
rect 423234 252308 423854 261398
rect 426954 265674 427574 272000
rect 428598 271829 428658 273670
rect 428595 271828 428661 271829
rect 428595 271764 428596 271828
rect 428660 271764 428661 271828
rect 428595 271763 428661 271764
rect 429702 270741 429762 273670
rect 430990 273325 431050 273670
rect 430987 273324 431053 273325
rect 430987 273260 430988 273324
rect 431052 273260 431053 273324
rect 430987 273259 431053 273260
rect 431174 271829 431234 273670
rect 432278 271829 432338 273670
rect 433382 271829 433442 273670
rect 433566 273670 433652 273730
rect 434408 273730 434468 274040
rect 435768 273730 435828 274040
rect 436040 273730 436100 274040
rect 436992 273730 437052 274040
rect 434408 273670 434730 273730
rect 435768 273670 435834 273730
rect 431171 271828 431237 271829
rect 431171 271764 431172 271828
rect 431236 271764 431237 271828
rect 431171 271763 431237 271764
rect 432275 271828 432341 271829
rect 432275 271764 432276 271828
rect 432340 271764 432341 271828
rect 432275 271763 432341 271764
rect 433379 271828 433445 271829
rect 433379 271764 433380 271828
rect 433444 271764 433445 271828
rect 433379 271763 433445 271764
rect 433566 271421 433626 273670
rect 433563 271420 433629 271421
rect 433563 271356 433564 271420
rect 433628 271356 433629 271420
rect 433563 271355 433629 271356
rect 429699 270740 429765 270741
rect 429699 270676 429700 270740
rect 429764 270676 429765 270740
rect 429699 270675 429765 270676
rect 426954 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 427574 265674
rect 426954 265354 427574 265438
rect 426954 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 427574 265354
rect 426954 252308 427574 265118
rect 433794 255454 434414 272000
rect 434670 270877 434730 273670
rect 434667 270876 434733 270877
rect 434667 270812 434668 270876
rect 434732 270812 434733 270876
rect 434667 270811 434733 270812
rect 435774 270741 435834 273670
rect 435958 273670 436100 273730
rect 436878 273670 437052 273730
rect 438080 273730 438140 274040
rect 438488 273730 438548 274040
rect 439168 273730 439228 274040
rect 440936 273730 440996 274040
rect 443520 273730 443580 274040
rect 438080 273670 438410 273730
rect 438488 273670 438594 273730
rect 439168 273670 439330 273730
rect 435958 271829 436018 273670
rect 435955 271828 436021 271829
rect 435955 271764 435956 271828
rect 436020 271764 436021 271828
rect 435955 271763 436021 271764
rect 436878 270877 436938 273670
rect 436875 270876 436941 270877
rect 436875 270812 436876 270876
rect 436940 270812 436941 270876
rect 436875 270811 436941 270812
rect 435771 270740 435837 270741
rect 435771 270676 435772 270740
rect 435836 270676 435837 270740
rect 435771 270675 435837 270676
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 252308 434414 254898
rect 437514 259174 438134 272000
rect 438350 270877 438410 273670
rect 438534 271829 438594 273670
rect 438531 271828 438597 271829
rect 438531 271764 438532 271828
rect 438596 271764 438597 271828
rect 438531 271763 438597 271764
rect 439270 271285 439330 273670
rect 440926 273670 440996 273730
rect 443502 273670 443580 273730
rect 440926 271421 440986 273670
rect 440923 271420 440989 271421
rect 440923 271356 440924 271420
rect 440988 271356 440989 271420
rect 440923 271355 440989 271356
rect 439267 271284 439333 271285
rect 439267 271220 439268 271284
rect 439332 271220 439333 271284
rect 439267 271219 439333 271220
rect 438347 270876 438413 270877
rect 438347 270812 438348 270876
rect 438412 270812 438413 270876
rect 438347 270811 438413 270812
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 252308 438134 258618
rect 441234 262894 441854 272000
rect 443502 271829 443562 273670
rect 445968 273597 446028 274040
rect 448280 273730 448340 274040
rect 451000 273730 451060 274040
rect 453448 273730 453508 274040
rect 455896 273730 455956 274040
rect 458480 273730 458540 274040
rect 448280 273670 448346 273730
rect 451000 273670 451106 273730
rect 445965 273596 446031 273597
rect 445965 273532 445966 273596
rect 446030 273532 446031 273596
rect 445965 273531 446031 273532
rect 443499 271828 443565 271829
rect 443499 271764 443500 271828
rect 443564 271764 443565 271828
rect 443499 271763 443565 271764
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 252308 441854 262338
rect 444954 266614 445574 272000
rect 448286 271829 448346 273670
rect 451046 271829 451106 273670
rect 453438 273670 453508 273730
rect 455830 273670 455956 273730
rect 458406 273670 458540 273730
rect 460928 273730 460988 274040
rect 463512 273730 463572 274040
rect 465960 273730 466020 274040
rect 468544 273730 468604 274040
rect 470992 273730 471052 274040
rect 460928 273670 461042 273730
rect 448283 271828 448349 271829
rect 448283 271764 448284 271828
rect 448348 271764 448349 271828
rect 448283 271763 448349 271764
rect 451043 271828 451109 271829
rect 451043 271764 451044 271828
rect 451108 271764 451109 271828
rect 451043 271763 451109 271764
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 252308 445574 266058
rect 451794 256394 452414 272000
rect 453438 271829 453498 273670
rect 455830 272237 455890 273670
rect 455827 272236 455893 272237
rect 455827 272172 455828 272236
rect 455892 272172 455893 272236
rect 455827 272171 455893 272172
rect 453435 271828 453501 271829
rect 453435 271764 453436 271828
rect 453500 271764 453501 271828
rect 453435 271763 453501 271764
rect 451794 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 452414 256394
rect 451794 256074 452414 256158
rect 451794 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 452414 256074
rect 451794 252308 452414 255838
rect 455514 260114 456134 272000
rect 458406 271829 458466 273670
rect 458403 271828 458469 271829
rect 458403 271764 458404 271828
rect 458468 271764 458469 271828
rect 458403 271763 458469 271764
rect 455514 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 456134 260114
rect 455514 259794 456134 259878
rect 455514 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 456134 259794
rect 455514 252308 456134 259558
rect 459234 261954 459854 272000
rect 460982 271557 461042 273670
rect 462638 273670 463572 273730
rect 465950 273670 466020 273730
rect 468526 273670 468604 273730
rect 470918 273670 471052 273730
rect 473440 273730 473500 274040
rect 475888 273730 475948 274040
rect 478472 273730 478532 274040
rect 480920 273730 480980 274040
rect 483368 273730 483428 274040
rect 473440 273670 473554 273730
rect 460979 271556 461045 271557
rect 460979 271492 460980 271556
rect 461044 271492 461045 271556
rect 460979 271491 461045 271492
rect 462638 271013 462698 273670
rect 462635 271012 462701 271013
rect 462635 270948 462636 271012
rect 462700 270948 462701 271012
rect 462635 270947 462701 270948
rect 459234 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 459854 261954
rect 459234 261634 459854 261718
rect 459234 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 459854 261634
rect 459234 252308 459854 261398
rect 462954 265674 463574 272000
rect 465950 271693 466010 273670
rect 468526 273053 468586 273670
rect 468523 273052 468589 273053
rect 468523 272988 468524 273052
rect 468588 272988 468589 273052
rect 468523 272987 468589 272988
rect 470918 272917 470978 273670
rect 470915 272916 470981 272917
rect 470915 272852 470916 272916
rect 470980 272852 470981 272916
rect 470915 272851 470981 272852
rect 473494 272781 473554 273670
rect 475886 273670 475948 273730
rect 478462 273670 478532 273730
rect 480854 273670 480980 273730
rect 483246 273670 483428 273730
rect 485952 273730 486012 274040
rect 503224 273730 503284 274040
rect 485952 273670 486066 273730
rect 473491 272780 473557 272781
rect 473491 272716 473492 272780
rect 473556 272716 473557 272780
rect 473491 272715 473557 272716
rect 475886 272645 475946 273670
rect 478462 272917 478522 273670
rect 478459 272916 478525 272917
rect 478459 272852 478460 272916
rect 478524 272852 478525 272916
rect 478459 272851 478525 272852
rect 480854 272781 480914 273670
rect 483246 273189 483306 273670
rect 483243 273188 483309 273189
rect 483243 273124 483244 273188
rect 483308 273124 483309 273188
rect 483243 273123 483309 273124
rect 480851 272780 480917 272781
rect 480851 272716 480852 272780
rect 480916 272716 480917 272780
rect 480851 272715 480917 272716
rect 486006 272645 486066 273670
rect 503118 273670 503284 273730
rect 503360 273730 503420 274040
rect 503360 273670 503546 273730
rect 475883 272644 475949 272645
rect 475883 272580 475884 272644
rect 475948 272580 475949 272644
rect 475883 272579 475949 272580
rect 486003 272644 486069 272645
rect 486003 272580 486004 272644
rect 486068 272580 486069 272644
rect 486003 272579 486069 272580
rect 465947 271692 466013 271693
rect 465947 271628 465948 271692
rect 466012 271628 466013 271692
rect 465947 271627 466013 271628
rect 462954 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 463574 265674
rect 462954 265354 463574 265438
rect 462954 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 463574 265354
rect 462954 252308 463574 265118
rect 469794 255454 470414 272000
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 252308 470414 254898
rect 473514 259174 474134 272000
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 252308 474134 258618
rect 477234 262894 477854 272000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 252308 477854 262338
rect 480954 266614 481574 272000
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 252308 481574 266058
rect 487794 256394 488414 272000
rect 487794 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 487794 256074 488414 256158
rect 487794 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 487794 252308 488414 255838
rect 491514 260114 492134 272000
rect 491514 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 491514 259794 492134 259878
rect 491514 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 491514 252308 492134 259558
rect 495234 261954 495854 272000
rect 495234 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 495234 261634 495854 261718
rect 495234 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 495234 252308 495854 261398
rect 498954 265674 499574 272000
rect 503118 271693 503178 273670
rect 503115 271692 503181 271693
rect 503115 271628 503116 271692
rect 503180 271628 503181 271692
rect 503115 271627 503181 271628
rect 503486 271285 503546 273670
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 503483 271284 503549 271285
rect 503483 271220 503484 271284
rect 503548 271220 503549 271284
rect 503483 271219 503549 271220
rect 498954 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 498954 265354 499574 265438
rect 498954 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 498515 252788 498581 252789
rect 498515 252724 498516 252788
rect 498580 252724 498581 252788
rect 498515 252723 498581 252724
rect 498518 250610 498578 252723
rect 498954 252308 499574 265118
rect 505794 255454 506414 272000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 499803 253332 499869 253333
rect 499803 253268 499804 253332
rect 499868 253268 499869 253332
rect 499803 253267 499869 253268
rect 499806 250610 499866 253267
rect 505794 252308 506414 254898
rect 509514 259174 510134 272000
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 252308 510134 258618
rect 513234 262894 513854 272000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 510843 252652 510909 252653
rect 510843 252588 510844 252652
rect 510908 252588 510909 252652
rect 510843 252587 510909 252588
rect 510846 250610 510906 252587
rect 513234 252308 513854 262338
rect 516954 266614 517574 272000
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 252308 517574 266058
rect 498464 250550 498578 250610
rect 499688 250550 499866 250610
rect 510840 250550 510906 250610
rect 498464 250240 498524 250550
rect 499688 250240 499748 250550
rect 510840 250240 510900 250550
rect 380272 237454 380620 237486
rect 380272 237218 380328 237454
rect 380564 237218 380620 237454
rect 380272 237134 380620 237218
rect 380272 236898 380328 237134
rect 380564 236898 380620 237134
rect 380272 236866 380620 236898
rect 516000 237454 516348 237486
rect 516000 237218 516056 237454
rect 516292 237218 516348 237454
rect 516000 237134 516348 237218
rect 516000 236898 516056 237134
rect 516292 236898 516348 237134
rect 516000 236866 516348 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 380952 219454 381300 219486
rect 380952 219218 381008 219454
rect 381244 219218 381300 219454
rect 380952 219134 381300 219218
rect 380952 218898 381008 219134
rect 381244 218898 381300 219134
rect 380952 218866 381300 218898
rect 515320 219454 515668 219486
rect 515320 219218 515376 219454
rect 515612 219218 515668 219454
rect 515320 219134 515668 219218
rect 515320 218898 515376 219134
rect 515612 218898 515668 219134
rect 515320 218866 515668 218898
rect 380272 201454 380620 201486
rect 380272 201218 380328 201454
rect 380564 201218 380620 201454
rect 380272 201134 380620 201218
rect 380272 200898 380328 201134
rect 380564 200898 380620 201134
rect 380272 200866 380620 200898
rect 516000 201454 516348 201486
rect 516000 201218 516056 201454
rect 516292 201218 516348 201454
rect 516000 201134 516348 201218
rect 516000 200898 516056 201134
rect 516292 200898 516348 201134
rect 516000 200866 516348 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 380952 183454 381300 183486
rect 380952 183218 381008 183454
rect 381244 183218 381300 183454
rect 380952 183134 381300 183218
rect 380952 182898 381008 183134
rect 381244 182898 381300 183134
rect 380952 182866 381300 182898
rect 515320 183454 515668 183486
rect 515320 183218 515376 183454
rect 515612 183218 515668 183454
rect 515320 183134 515668 183218
rect 515320 182898 515376 183134
rect 515612 182898 515668 183134
rect 515320 182866 515668 182898
rect 379470 171090 379714 171150
rect 379470 165069 379530 171090
rect 396056 167010 396116 167106
rect 397144 167010 397204 167106
rect 396030 166950 396116 167010
rect 397134 166950 397204 167010
rect 398232 167010 398292 167106
rect 399592 167010 399652 167106
rect 400544 167010 400604 167106
rect 401768 167010 401828 167106
rect 403128 167010 403188 167106
rect 404216 167010 404276 167106
rect 405440 167010 405500 167106
rect 406528 167010 406588 167106
rect 398232 166950 398298 167010
rect 379467 165068 379533 165069
rect 379467 165004 379468 165068
rect 379532 165004 379533 165068
rect 379467 165003 379533 165004
rect 379794 148394 380414 165000
rect 379794 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 380414 148394
rect 379794 148074 380414 148158
rect 379794 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 380414 148074
rect 379467 146164 379533 146165
rect 379467 146100 379468 146164
rect 379532 146100 379533 146164
rect 379467 146099 379533 146100
rect 379470 145621 379530 146099
rect 379467 145620 379533 145621
rect 379467 145556 379468 145620
rect 379532 145556 379533 145620
rect 379467 145555 379533 145556
rect 379470 142170 379530 145555
rect 379794 145308 380414 147838
rect 383514 152114 384134 165000
rect 383514 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 384134 152114
rect 383514 151794 384134 151878
rect 383514 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 384134 151794
rect 383514 145308 384134 151558
rect 387234 155834 387854 165000
rect 387234 155598 387266 155834
rect 387502 155598 387586 155834
rect 387822 155598 387854 155834
rect 387234 155514 387854 155598
rect 387234 155278 387266 155514
rect 387502 155278 387586 155514
rect 387822 155278 387854 155514
rect 387234 145308 387854 155278
rect 390954 157674 391574 165000
rect 396030 164253 396090 166950
rect 397134 164389 397194 166950
rect 398238 165613 398298 166950
rect 399526 166950 399652 167010
rect 400446 166950 400604 167010
rect 401734 166950 401828 167010
rect 403022 166950 403188 167010
rect 404126 166950 404276 167010
rect 405414 166950 405500 167010
rect 406518 166950 406588 167010
rect 407616 167010 407676 167106
rect 408296 167010 408356 167106
rect 407616 166950 407682 167010
rect 398235 165612 398301 165613
rect 398235 165548 398236 165612
rect 398300 165548 398301 165612
rect 398235 165547 398301 165548
rect 397131 164388 397197 164389
rect 397131 164324 397132 164388
rect 397196 164324 397197 164388
rect 397131 164323 397197 164324
rect 396027 164252 396093 164253
rect 396027 164188 396028 164252
rect 396092 164188 396093 164252
rect 396027 164187 396093 164188
rect 390954 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 391574 157674
rect 390954 157354 391574 157438
rect 390954 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 391574 157354
rect 390954 145308 391574 157118
rect 397794 147454 398414 165000
rect 399526 164253 399586 166950
rect 400446 164253 400506 166950
rect 401734 165613 401794 166950
rect 401731 165612 401797 165613
rect 401731 165548 401732 165612
rect 401796 165548 401797 165612
rect 401731 165547 401797 165548
rect 399523 164252 399589 164253
rect 399523 164188 399524 164252
rect 399588 164188 399589 164252
rect 399523 164187 399589 164188
rect 400443 164252 400509 164253
rect 400443 164188 400444 164252
rect 400508 164188 400509 164252
rect 400443 164187 400509 164188
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 145308 398414 146898
rect 401514 151174 402134 165000
rect 403022 164253 403082 166950
rect 404126 164389 404186 166950
rect 405414 165613 405474 166950
rect 405411 165612 405477 165613
rect 405411 165548 405412 165612
rect 405476 165548 405477 165612
rect 405411 165547 405477 165548
rect 404123 164388 404189 164389
rect 404123 164324 404124 164388
rect 404188 164324 404189 164388
rect 404123 164323 404189 164324
rect 403019 164252 403085 164253
rect 403019 164188 403020 164252
rect 403084 164188 403085 164252
rect 403019 164187 403085 164188
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 145308 402134 150618
rect 405234 154894 405854 165000
rect 406518 164253 406578 166950
rect 407622 164253 407682 166950
rect 408174 166950 408356 167010
rect 408704 167010 408764 167106
rect 410064 167010 410124 167106
rect 408704 166950 408786 167010
rect 408174 165613 408234 166950
rect 408171 165612 408237 165613
rect 408171 165548 408172 165612
rect 408236 165548 408237 165612
rect 408171 165547 408237 165548
rect 408726 164253 408786 166950
rect 410014 166950 410124 167010
rect 410744 167010 410804 167106
rect 411288 167010 411348 167106
rect 412376 167010 412436 167106
rect 413464 167010 413524 167106
rect 410744 166950 410810 167010
rect 411288 166950 411362 167010
rect 412376 166950 412466 167010
rect 406515 164252 406581 164253
rect 406515 164188 406516 164252
rect 406580 164188 406581 164252
rect 406515 164187 406581 164188
rect 407619 164252 407685 164253
rect 407619 164188 407620 164252
rect 407684 164188 407685 164252
rect 407619 164187 407685 164188
rect 408723 164252 408789 164253
rect 408723 164188 408724 164252
rect 408788 164188 408789 164252
rect 408723 164187 408789 164188
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 145308 405854 154338
rect 408954 158614 409574 165000
rect 410014 164253 410074 166950
rect 410750 164797 410810 166950
rect 410747 164796 410813 164797
rect 410747 164732 410748 164796
rect 410812 164732 410813 164796
rect 410747 164731 410813 164732
rect 411302 164253 411362 166950
rect 412406 164389 412466 166950
rect 413326 166950 413524 167010
rect 413600 167010 413660 167106
rect 414552 167010 414612 167106
rect 415912 167010 415972 167106
rect 413600 166950 413754 167010
rect 412403 164388 412469 164389
rect 412403 164324 412404 164388
rect 412468 164324 412469 164388
rect 412403 164323 412469 164324
rect 413326 164253 413386 166950
rect 413694 164933 413754 166950
rect 414430 166950 414612 167010
rect 415902 166950 415972 167010
rect 416048 167010 416108 167106
rect 417000 167010 417060 167106
rect 418088 167010 418148 167106
rect 418496 167010 418556 167106
rect 419448 167010 419508 167106
rect 416048 166950 416146 167010
rect 417000 166950 417066 167010
rect 418088 166950 418354 167010
rect 413691 164932 413757 164933
rect 413691 164868 413692 164932
rect 413756 164868 413757 164932
rect 413691 164867 413757 164868
rect 414430 164253 414490 166950
rect 415902 165613 415962 166950
rect 416086 165613 416146 166950
rect 415899 165612 415965 165613
rect 415899 165548 415900 165612
rect 415964 165548 415965 165612
rect 415899 165547 415965 165548
rect 416083 165612 416149 165613
rect 416083 165548 416084 165612
rect 416148 165548 416149 165612
rect 416083 165547 416149 165548
rect 410011 164252 410077 164253
rect 410011 164188 410012 164252
rect 410076 164188 410077 164252
rect 410011 164187 410077 164188
rect 411299 164252 411365 164253
rect 411299 164188 411300 164252
rect 411364 164188 411365 164252
rect 411299 164187 411365 164188
rect 413323 164252 413389 164253
rect 413323 164188 413324 164252
rect 413388 164188 413389 164252
rect 413323 164187 413389 164188
rect 414427 164252 414493 164253
rect 414427 164188 414428 164252
rect 414492 164188 414493 164252
rect 414427 164187 414493 164188
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 145308 409574 158058
rect 415794 148394 416414 165000
rect 417006 164253 417066 166950
rect 418294 164253 418354 166950
rect 418478 166950 418556 167010
rect 419398 166950 419508 167010
rect 420672 167010 420732 167106
rect 421080 167010 421140 167106
rect 420672 166950 420746 167010
rect 418478 166837 418538 166950
rect 418475 166836 418541 166837
rect 418475 166772 418476 166836
rect 418540 166772 418541 166836
rect 418475 166771 418541 166772
rect 419398 165613 419458 166950
rect 419395 165612 419461 165613
rect 419395 165548 419396 165612
rect 419460 165548 419461 165612
rect 419395 165547 419461 165548
rect 417003 164252 417069 164253
rect 417003 164188 417004 164252
rect 417068 164188 417069 164252
rect 417003 164187 417069 164188
rect 418291 164252 418357 164253
rect 418291 164188 418292 164252
rect 418356 164188 418357 164252
rect 418291 164187 418357 164188
rect 415794 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 416414 148394
rect 415794 148074 416414 148158
rect 415794 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 416414 148074
rect 415794 145308 416414 147838
rect 419514 152114 420134 165000
rect 420686 164253 420746 166950
rect 421054 166950 421140 167010
rect 421760 167010 421820 167106
rect 422848 167010 422908 167106
rect 423528 167010 423588 167106
rect 423936 167010 423996 167106
rect 425296 167010 425356 167106
rect 421760 166950 421850 167010
rect 422848 166950 422954 167010
rect 421054 166837 421114 166950
rect 421051 166836 421117 166837
rect 421051 166772 421052 166836
rect 421116 166772 421117 166836
rect 421051 166771 421117 166772
rect 421790 164525 421850 166950
rect 421787 164524 421853 164525
rect 421787 164460 421788 164524
rect 421852 164460 421853 164524
rect 421787 164459 421853 164460
rect 422894 164253 422954 166950
rect 423446 166950 423588 167010
rect 423814 166950 423996 167010
rect 425286 166950 425356 167010
rect 425976 167010 426036 167106
rect 426384 167010 426444 167106
rect 427608 167010 427668 167106
rect 425976 166950 426082 167010
rect 426384 166950 426450 167010
rect 423446 166293 423506 166950
rect 423443 166292 423509 166293
rect 423443 166228 423444 166292
rect 423508 166228 423509 166292
rect 423443 166227 423509 166228
rect 423814 165613 423874 166950
rect 423811 165612 423877 165613
rect 423811 165548 423812 165612
rect 423876 165548 423877 165612
rect 423811 165547 423877 165548
rect 420683 164252 420749 164253
rect 420683 164188 420684 164252
rect 420748 164188 420749 164252
rect 420683 164187 420749 164188
rect 422891 164252 422957 164253
rect 422891 164188 422892 164252
rect 422956 164188 422957 164252
rect 422891 164187 422957 164188
rect 419514 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 420134 152114
rect 419514 151794 420134 151878
rect 419514 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 420134 151794
rect 419514 145308 420134 151558
rect 423234 155834 423854 165000
rect 425286 164253 425346 166950
rect 426022 165069 426082 166950
rect 426019 165068 426085 165069
rect 426019 165004 426020 165068
rect 426084 165004 426085 165068
rect 426019 165003 426085 165004
rect 426390 164253 426450 166950
rect 427494 166950 427668 167010
rect 427494 165613 427554 166950
rect 428288 166837 428348 167106
rect 428285 166836 428351 166837
rect 428285 166772 428286 166836
rect 428350 166772 428351 166836
rect 428285 166771 428351 166772
rect 428696 166290 428756 167106
rect 429784 166290 429844 167106
rect 431008 166837 431068 167106
rect 431005 166836 431071 166837
rect 431005 166772 431006 166836
rect 431070 166772 431071 166836
rect 431005 166771 431071 166772
rect 428696 166230 428842 166290
rect 427491 165612 427557 165613
rect 427491 165548 427492 165612
rect 427556 165548 427557 165612
rect 427491 165547 427557 165548
rect 425283 164252 425349 164253
rect 425283 164188 425284 164252
rect 425348 164188 425349 164252
rect 425283 164187 425349 164188
rect 426387 164252 426453 164253
rect 426387 164188 426388 164252
rect 426452 164188 426453 164252
rect 426387 164187 426453 164188
rect 423234 155598 423266 155834
rect 423502 155598 423586 155834
rect 423822 155598 423854 155834
rect 423234 155514 423854 155598
rect 423234 155278 423266 155514
rect 423502 155278 423586 155514
rect 423822 155278 423854 155514
rect 423234 145308 423854 155278
rect 426954 157674 427574 165000
rect 428782 164253 428842 166230
rect 429702 166230 429844 166290
rect 431144 166290 431204 167106
rect 432232 166290 432292 167106
rect 433320 166290 433380 167106
rect 433592 166837 433652 167106
rect 433589 166836 433655 166837
rect 433589 166772 433590 166836
rect 433654 166772 433655 166836
rect 433589 166771 433655 166772
rect 434408 166565 434468 167106
rect 434405 166564 434471 166565
rect 434405 166500 434406 166564
rect 434470 166500 434471 166564
rect 434405 166499 434471 166500
rect 435768 166290 435828 167106
rect 436040 166290 436100 167106
rect 436992 166290 437052 167106
rect 438080 166290 438140 167106
rect 431144 166230 431234 166290
rect 432232 166230 432338 166290
rect 433320 166230 433442 166290
rect 435768 166230 435834 166290
rect 429702 165613 429762 166230
rect 429699 165612 429765 165613
rect 429699 165548 429700 165612
rect 429764 165548 429765 165612
rect 429699 165547 429765 165548
rect 431174 164525 431234 166230
rect 432278 165069 432338 166230
rect 432275 165068 432341 165069
rect 432275 165004 432276 165068
rect 432340 165004 432341 165068
rect 432275 165003 432341 165004
rect 431171 164524 431237 164525
rect 431171 164460 431172 164524
rect 431236 164460 431237 164524
rect 431171 164459 431237 164460
rect 433382 164253 433442 166230
rect 435774 165613 435834 166230
rect 435958 166230 436100 166290
rect 436878 166230 437052 166290
rect 437982 166230 438140 166290
rect 438488 166290 438548 167106
rect 439168 166290 439228 167106
rect 440936 166290 440996 167106
rect 443520 166290 443580 167106
rect 445968 166290 446028 167106
rect 448280 167010 448340 167106
rect 451000 167010 451060 167106
rect 453448 167010 453508 167106
rect 455896 167010 455956 167106
rect 448280 166950 448346 167010
rect 451000 166950 451106 167010
rect 438488 166230 438594 166290
rect 439168 166230 439330 166290
rect 435958 165613 436018 166230
rect 435771 165612 435837 165613
rect 435771 165548 435772 165612
rect 435836 165548 435837 165612
rect 435771 165547 435837 165548
rect 435955 165612 436021 165613
rect 435955 165548 435956 165612
rect 436020 165548 436021 165612
rect 435955 165547 436021 165548
rect 428779 164252 428845 164253
rect 428779 164188 428780 164252
rect 428844 164188 428845 164252
rect 428779 164187 428845 164188
rect 433379 164252 433445 164253
rect 433379 164188 433380 164252
rect 433444 164188 433445 164252
rect 433379 164187 433445 164188
rect 426954 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 427574 157674
rect 426954 157354 427574 157438
rect 426954 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 427574 157354
rect 426954 145308 427574 157118
rect 433794 147454 434414 165000
rect 436878 164933 436938 166230
rect 437982 165613 438042 166230
rect 438534 165613 438594 166230
rect 439270 165613 439330 166230
rect 440926 166230 440996 166290
rect 443502 166230 443580 166290
rect 445894 166230 446028 166290
rect 440926 165613 440986 166230
rect 443502 165613 443562 166230
rect 445894 165613 445954 166230
rect 448286 165613 448346 166950
rect 451046 165613 451106 166950
rect 453438 166950 453508 167010
rect 455830 166950 455956 167010
rect 453438 165613 453498 166950
rect 455830 165613 455890 166950
rect 458480 166290 458540 167106
rect 458406 166230 458540 166290
rect 460928 166290 460988 167106
rect 463512 166290 463572 167106
rect 465960 166290 466020 167106
rect 468544 166290 468604 167106
rect 470992 166837 471052 167106
rect 473440 166837 473500 167106
rect 475888 166837 475948 167106
rect 478472 166837 478532 167106
rect 480920 166837 480980 167106
rect 470989 166836 471055 166837
rect 470989 166772 470990 166836
rect 471054 166772 471055 166836
rect 470989 166771 471055 166772
rect 473437 166836 473503 166837
rect 473437 166772 473438 166836
rect 473502 166772 473503 166836
rect 473437 166771 473503 166772
rect 475885 166836 475951 166837
rect 475885 166772 475886 166836
rect 475950 166772 475951 166836
rect 475885 166771 475951 166772
rect 478469 166836 478535 166837
rect 478469 166772 478470 166836
rect 478534 166772 478535 166836
rect 478469 166771 478535 166772
rect 480917 166836 480983 166837
rect 480917 166772 480918 166836
rect 480982 166772 480983 166836
rect 480917 166771 480983 166772
rect 483368 166701 483428 167106
rect 485952 166701 486012 167106
rect 483365 166700 483431 166701
rect 483365 166636 483366 166700
rect 483430 166636 483431 166700
rect 483365 166635 483431 166636
rect 485949 166700 486015 166701
rect 485949 166636 485950 166700
rect 486014 166636 486015 166700
rect 485949 166635 486015 166636
rect 503224 166565 503284 167106
rect 503221 166564 503287 166565
rect 503221 166500 503222 166564
rect 503286 166500 503287 166564
rect 503221 166499 503287 166500
rect 503360 166290 503420 167106
rect 460928 166230 461042 166290
rect 463512 166230 463618 166290
rect 458406 165613 458466 166230
rect 437979 165612 438045 165613
rect 437979 165548 437980 165612
rect 438044 165548 438045 165612
rect 437979 165547 438045 165548
rect 438531 165612 438597 165613
rect 438531 165548 438532 165612
rect 438596 165548 438597 165612
rect 438531 165547 438597 165548
rect 439267 165612 439333 165613
rect 439267 165548 439268 165612
rect 439332 165548 439333 165612
rect 439267 165547 439333 165548
rect 440923 165612 440989 165613
rect 440923 165548 440924 165612
rect 440988 165548 440989 165612
rect 440923 165547 440989 165548
rect 443499 165612 443565 165613
rect 443499 165548 443500 165612
rect 443564 165548 443565 165612
rect 443499 165547 443565 165548
rect 445891 165612 445957 165613
rect 445891 165548 445892 165612
rect 445956 165548 445957 165612
rect 445891 165547 445957 165548
rect 448283 165612 448349 165613
rect 448283 165548 448284 165612
rect 448348 165548 448349 165612
rect 448283 165547 448349 165548
rect 451043 165612 451109 165613
rect 451043 165548 451044 165612
rect 451108 165548 451109 165612
rect 451043 165547 451109 165548
rect 453435 165612 453501 165613
rect 453435 165548 453436 165612
rect 453500 165548 453501 165612
rect 453435 165547 453501 165548
rect 455827 165612 455893 165613
rect 455827 165548 455828 165612
rect 455892 165548 455893 165612
rect 455827 165547 455893 165548
rect 458403 165612 458469 165613
rect 458403 165548 458404 165612
rect 458468 165548 458469 165612
rect 458403 165547 458469 165548
rect 436875 164932 436941 164933
rect 436875 164868 436876 164932
rect 436940 164868 436941 164932
rect 436875 164867 436941 164868
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 145308 434414 146898
rect 437514 151174 438134 165000
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 145308 438134 150618
rect 441234 154894 441854 165000
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 145308 441854 154338
rect 444954 158614 445574 165000
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 145308 445574 158058
rect 451794 148394 452414 165000
rect 451794 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 452414 148394
rect 451794 148074 452414 148158
rect 451794 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 452414 148074
rect 451794 145308 452414 147838
rect 455514 152114 456134 165000
rect 455514 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 456134 152114
rect 455514 151794 456134 151878
rect 455514 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 456134 151794
rect 455514 145308 456134 151558
rect 459234 155834 459854 165000
rect 460982 164661 461042 166230
rect 463558 165205 463618 166230
rect 465950 166230 466020 166290
rect 468526 166230 468604 166290
rect 503302 166230 503420 166290
rect 465950 165341 466010 166230
rect 468526 165477 468586 166230
rect 503302 165613 503362 166230
rect 503299 165612 503365 165613
rect 503299 165548 503300 165612
rect 503364 165548 503365 165612
rect 503299 165547 503365 165548
rect 468523 165476 468589 165477
rect 468523 165412 468524 165476
rect 468588 165412 468589 165476
rect 468523 165411 468589 165412
rect 523794 165454 524414 200898
rect 465947 165340 466013 165341
rect 465947 165276 465948 165340
rect 466012 165276 466013 165340
rect 465947 165275 466013 165276
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 463555 165204 463621 165205
rect 463555 165140 463556 165204
rect 463620 165140 463621 165204
rect 463555 165139 463621 165140
rect 523794 165134 524414 165218
rect 460979 164660 461045 164661
rect 460979 164596 460980 164660
rect 461044 164596 461045 164660
rect 460979 164595 461045 164596
rect 459234 155598 459266 155834
rect 459502 155598 459586 155834
rect 459822 155598 459854 155834
rect 459234 155514 459854 155598
rect 459234 155278 459266 155514
rect 459502 155278 459586 155514
rect 459822 155278 459854 155514
rect 459234 145308 459854 155278
rect 462954 157674 463574 165000
rect 462954 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 463574 157674
rect 462954 157354 463574 157438
rect 462954 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 463574 157354
rect 462954 145308 463574 157118
rect 469794 147454 470414 165000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 145308 470414 146898
rect 473514 151174 474134 165000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 145308 474134 150618
rect 477234 154894 477854 165000
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 145308 477854 154338
rect 480954 158614 481574 165000
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 145308 481574 158058
rect 487794 148394 488414 165000
rect 487794 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 487794 148074 488414 148158
rect 487794 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 487794 145308 488414 147838
rect 491514 152114 492134 165000
rect 491514 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 491514 151794 492134 151878
rect 491514 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 491514 145308 492134 151558
rect 495234 155834 495854 165000
rect 495234 155598 495266 155834
rect 495502 155598 495586 155834
rect 495822 155598 495854 155834
rect 495234 155514 495854 155598
rect 495234 155278 495266 155514
rect 495502 155278 495586 155514
rect 495822 155278 495854 155514
rect 495234 145308 495854 155278
rect 498954 157674 499574 165000
rect 498954 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 498954 157354 499574 157438
rect 498954 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 498954 145308 499574 157118
rect 505794 147454 506414 165000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 145308 506414 146898
rect 509514 151174 510134 165000
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 145308 510134 150618
rect 513234 154894 513854 165000
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 510843 145484 510909 145485
rect 510843 145420 510844 145484
rect 510908 145420 510909 145484
rect 510843 145419 510909 145420
rect 498515 144940 498581 144941
rect 498515 144876 498516 144940
rect 498580 144876 498581 144940
rect 498515 144875 498581 144876
rect 499803 144940 499869 144941
rect 499803 144876 499804 144940
rect 499868 144876 499869 144940
rect 499803 144875 499869 144876
rect 498518 143850 498578 144875
rect 499806 143850 499866 144875
rect 510846 143850 510906 145419
rect 513234 145308 513854 154338
rect 516954 158614 517574 165000
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 145308 517574 158058
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 498464 143790 498578 143850
rect 499688 143790 499866 143850
rect 510840 143790 510906 143850
rect 498464 143202 498524 143790
rect 499688 143202 499748 143790
rect 510840 143202 510900 143790
rect 379470 142110 379714 142170
rect 379654 64890 379714 142110
rect 380272 129454 380620 129486
rect 380272 129218 380328 129454
rect 380564 129218 380620 129454
rect 380272 129134 380620 129218
rect 380272 128898 380328 129134
rect 380564 128898 380620 129134
rect 380272 128866 380620 128898
rect 516000 129454 516348 129486
rect 516000 129218 516056 129454
rect 516292 129218 516348 129454
rect 516000 129134 516348 129218
rect 516000 128898 516056 129134
rect 516292 128898 516348 129134
rect 516000 128866 516348 128898
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 380952 111454 381300 111486
rect 380952 111218 381008 111454
rect 381244 111218 381300 111454
rect 380952 111134 381300 111218
rect 380952 110898 381008 111134
rect 381244 110898 381300 111134
rect 380952 110866 381300 110898
rect 515320 111454 515668 111486
rect 515320 111218 515376 111454
rect 515612 111218 515668 111454
rect 515320 111134 515668 111218
rect 515320 110898 515376 111134
rect 515612 110898 515668 111134
rect 515320 110866 515668 110898
rect 380272 93454 380620 93486
rect 380272 93218 380328 93454
rect 380564 93218 380620 93454
rect 380272 93134 380620 93218
rect 380272 92898 380328 93134
rect 380564 92898 380620 93134
rect 380272 92866 380620 92898
rect 516000 93454 516348 93486
rect 516000 93218 516056 93454
rect 516292 93218 516348 93454
rect 516000 93134 516348 93218
rect 516000 92898 516056 93134
rect 516292 92898 516348 93134
rect 516000 92866 516348 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 380952 75454 381300 75486
rect 380952 75218 381008 75454
rect 381244 75218 381300 75454
rect 380952 75134 381300 75218
rect 380952 74898 381008 75134
rect 381244 74898 381300 75134
rect 380952 74866 381300 74898
rect 515320 75454 515668 75486
rect 515320 75218 515376 75454
rect 515612 75218 515668 75454
rect 515320 75134 515668 75218
rect 515320 74898 515376 75134
rect 515612 74898 515668 75134
rect 515320 74866 515668 74898
rect 379470 64830 379714 64890
rect 379099 57356 379165 57357
rect 379099 57292 379100 57356
rect 379164 57292 379165 57356
rect 379099 57291 379165 57292
rect 378915 57220 378981 57221
rect 378915 57156 378916 57220
rect 378980 57156 378981 57220
rect 378915 57155 378981 57156
rect 378731 57084 378797 57085
rect 378731 57020 378732 57084
rect 378796 57020 378797 57084
rect 378731 57019 378797 57020
rect 379470 56133 379530 64830
rect 396056 59805 396116 60106
rect 397144 59805 397204 60106
rect 396053 59804 396119 59805
rect 396053 59740 396054 59804
rect 396118 59740 396119 59804
rect 396053 59739 396119 59740
rect 397141 59804 397207 59805
rect 397141 59740 397142 59804
rect 397206 59740 397207 59804
rect 397141 59739 397207 59740
rect 398232 59530 398292 60106
rect 399592 59802 399652 60106
rect 400544 59802 400604 60106
rect 399526 59742 399652 59802
rect 400446 59742 400604 59802
rect 398232 59470 398298 59530
rect 398238 58173 398298 59470
rect 398235 58172 398301 58173
rect 398235 58108 398236 58172
rect 398300 58108 398301 58172
rect 398235 58107 398301 58108
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379467 56132 379533 56133
rect 379467 56068 379468 56132
rect 379532 56068 379533 56132
rect 379467 56067 379533 56068
rect 377811 55996 377877 55997
rect 377811 55932 377812 55996
rect 377876 55932 377877 55996
rect 377811 55931 377877 55932
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 399526 57901 399586 59742
rect 400446 57901 400506 59742
rect 401768 59530 401828 60106
rect 403128 59805 403188 60106
rect 403125 59804 403191 59805
rect 403125 59740 403126 59804
rect 403190 59740 403191 59804
rect 403125 59739 403191 59740
rect 404216 59669 404276 60106
rect 404213 59668 404279 59669
rect 404213 59604 404214 59668
rect 404278 59604 404279 59668
rect 404213 59603 404279 59604
rect 405440 59530 405500 60106
rect 406528 59530 406588 60106
rect 401734 59470 401828 59530
rect 405414 59470 405500 59530
rect 406518 59470 406588 59530
rect 407616 59530 407676 60106
rect 408296 59530 408356 60106
rect 408704 59530 408764 60106
rect 410064 59530 410124 60106
rect 407616 59470 407682 59530
rect 408296 59470 408418 59530
rect 408704 59470 408786 59530
rect 401734 58173 401794 59470
rect 405414 58173 405474 59470
rect 401731 58172 401797 58173
rect 401731 58108 401732 58172
rect 401796 58108 401797 58172
rect 401731 58107 401797 58108
rect 405411 58172 405477 58173
rect 405411 58108 405412 58172
rect 405476 58108 405477 58172
rect 405411 58107 405477 58108
rect 399523 57900 399589 57901
rect 399523 57836 399524 57900
rect 399588 57836 399589 57900
rect 399523 57835 399589 57836
rect 400443 57900 400509 57901
rect 400443 57836 400444 57900
rect 400508 57836 400509 57900
rect 400443 57835 400509 57836
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 406518 57901 406578 59470
rect 407622 57901 407682 59470
rect 408358 57901 408418 59470
rect 408726 57901 408786 59470
rect 410014 59470 410124 59530
rect 410744 59530 410804 60106
rect 411288 59530 411348 60106
rect 412376 59530 412436 60106
rect 413464 59669 413524 60106
rect 413461 59668 413527 59669
rect 413461 59604 413462 59668
rect 413526 59604 413527 59668
rect 413461 59603 413527 59604
rect 413600 59530 413660 60106
rect 410744 59470 410810 59530
rect 411288 59470 411362 59530
rect 412376 59470 412466 59530
rect 406515 57900 406581 57901
rect 406515 57836 406516 57900
rect 406580 57836 406581 57900
rect 406515 57835 406581 57836
rect 407619 57900 407685 57901
rect 407619 57836 407620 57900
rect 407684 57836 407685 57900
rect 407619 57835 407685 57836
rect 408355 57900 408421 57901
rect 408355 57836 408356 57900
rect 408420 57836 408421 57900
rect 408355 57835 408421 57836
rect 408723 57900 408789 57901
rect 408723 57836 408724 57900
rect 408788 57836 408789 57900
rect 408723 57835 408789 57836
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 410014 57901 410074 59470
rect 410750 59397 410810 59470
rect 410747 59396 410813 59397
rect 410747 59332 410748 59396
rect 410812 59332 410813 59396
rect 410747 59331 410813 59332
rect 410011 57900 410077 57901
rect 410011 57836 410012 57900
rect 410076 57836 410077 57900
rect 410011 57835 410077 57836
rect 411302 56949 411362 59470
rect 412406 57901 412466 59470
rect 413510 59470 413660 59530
rect 414552 59530 414612 60106
rect 415912 59530 415972 60106
rect 414552 59470 414674 59530
rect 412403 57900 412469 57901
rect 412403 57836 412404 57900
rect 412468 57836 412469 57900
rect 412403 57835 412469 57836
rect 413510 57085 413570 59470
rect 414614 59397 414674 59470
rect 415534 59470 415972 59530
rect 416048 59530 416108 60106
rect 417000 59805 417060 60106
rect 416997 59804 417063 59805
rect 416997 59740 416998 59804
rect 417062 59740 417063 59804
rect 416997 59739 417063 59740
rect 418088 59530 418148 60106
rect 418496 59530 418556 60106
rect 419448 59530 419508 60106
rect 416048 59470 416146 59530
rect 418088 59470 418170 59530
rect 414611 59396 414677 59397
rect 414611 59332 414612 59396
rect 414676 59332 414677 59396
rect 414611 59331 414677 59332
rect 415534 57901 415594 59470
rect 416086 59397 416146 59470
rect 418110 59397 418170 59470
rect 418478 59470 418556 59530
rect 419398 59470 419508 59530
rect 420672 59530 420732 60106
rect 421080 59530 421140 60106
rect 420672 59470 420746 59530
rect 416083 59396 416149 59397
rect 416083 59332 416084 59396
rect 416148 59332 416149 59396
rect 416083 59331 416149 59332
rect 418107 59396 418173 59397
rect 418107 59332 418108 59396
rect 418172 59332 418173 59396
rect 418107 59331 418173 59332
rect 415531 57900 415597 57901
rect 415531 57836 415532 57900
rect 415596 57836 415597 57900
rect 415531 57835 415597 57836
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 418478 57221 418538 59470
rect 419398 59397 419458 59470
rect 420686 59397 420746 59470
rect 421054 59470 421140 59530
rect 421760 59530 421820 60106
rect 422848 59805 422908 60106
rect 422845 59804 422911 59805
rect 422845 59740 422846 59804
rect 422910 59740 422911 59804
rect 422845 59739 422911 59740
rect 423528 59669 423588 60106
rect 423936 59805 423996 60106
rect 423933 59804 423999 59805
rect 423933 59740 423934 59804
rect 423998 59740 423999 59804
rect 423933 59739 423999 59740
rect 423525 59668 423591 59669
rect 423525 59604 423526 59668
rect 423590 59604 423591 59668
rect 423525 59603 423591 59604
rect 425296 59530 425356 60106
rect 421760 59470 421850 59530
rect 419395 59396 419461 59397
rect 419395 59332 419396 59396
rect 419460 59332 419461 59396
rect 419395 59331 419461 59332
rect 420683 59396 420749 59397
rect 420683 59332 420684 59396
rect 420748 59332 420749 59396
rect 420683 59331 420749 59332
rect 415794 57134 416414 57218
rect 418475 57220 418541 57221
rect 418475 57156 418476 57220
rect 418540 57156 418541 57220
rect 418475 57155 418541 57156
rect 413507 57084 413573 57085
rect 413507 57020 413508 57084
rect 413572 57020 413573 57084
rect 413507 57019 413573 57020
rect 411299 56948 411365 56949
rect 411299 56884 411300 56948
rect 411364 56884 411365 56948
rect 411299 56883 411365 56884
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 421054 56405 421114 59470
rect 421790 59397 421850 59470
rect 425286 59470 425356 59530
rect 425976 59530 426036 60106
rect 426384 59530 426444 60106
rect 427608 59530 427668 60106
rect 428288 59530 428348 60106
rect 428696 59530 428756 60106
rect 429784 59530 429844 60106
rect 431008 59530 431068 60106
rect 425976 59470 426082 59530
rect 426384 59470 426450 59530
rect 427608 59470 427738 59530
rect 421787 59396 421853 59397
rect 421787 59332 421788 59396
rect 421852 59332 421853 59396
rect 421787 59331 421853 59332
rect 421051 56404 421117 56405
rect 421051 56340 421052 56404
rect 421116 56340 421117 56404
rect 421051 56339 421117 56340
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 425286 57901 425346 59470
rect 425283 57900 425349 57901
rect 425283 57836 425284 57900
rect 425348 57836 425349 57900
rect 425283 57835 425349 57836
rect 426022 56541 426082 59470
rect 426390 57901 426450 59470
rect 426387 57900 426453 57901
rect 426387 57836 426388 57900
rect 426452 57836 426453 57900
rect 426387 57835 426453 57836
rect 426019 56540 426085 56541
rect 426019 56476 426020 56540
rect 426084 56476 426085 56540
rect 426019 56475 426085 56476
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 427678 57221 427738 59470
rect 428230 59470 428348 59530
rect 428598 59470 428756 59530
rect 429702 59470 429844 59530
rect 430990 59470 431068 59530
rect 431144 59530 431204 60106
rect 432232 59530 432292 60106
rect 433320 59530 433380 60106
rect 433592 59530 433652 60106
rect 431144 59470 431234 59530
rect 432232 59470 432338 59530
rect 433320 59470 433442 59530
rect 428230 59397 428290 59470
rect 428227 59396 428293 59397
rect 428227 59332 428228 59396
rect 428292 59332 428293 59396
rect 428227 59331 428293 59332
rect 428598 57901 428658 59470
rect 429702 57901 429762 59470
rect 428595 57900 428661 57901
rect 428595 57836 428596 57900
rect 428660 57836 428661 57900
rect 428595 57835 428661 57836
rect 429699 57900 429765 57901
rect 429699 57836 429700 57900
rect 429764 57836 429765 57900
rect 429699 57835 429765 57836
rect 430990 57221 431050 59470
rect 431174 57901 431234 59470
rect 432278 57901 432338 59470
rect 431171 57900 431237 57901
rect 431171 57836 431172 57900
rect 431236 57836 431237 57900
rect 431171 57835 431237 57836
rect 432275 57900 432341 57901
rect 432275 57836 432276 57900
rect 432340 57836 432341 57900
rect 432275 57835 432341 57836
rect 433382 57493 433442 59470
rect 433566 59470 433652 59530
rect 434408 59530 434468 60106
rect 435768 59530 435828 60106
rect 436040 59530 436100 60106
rect 436992 59530 437052 60106
rect 434408 59470 434730 59530
rect 435768 59470 435834 59530
rect 433566 57901 433626 59470
rect 433563 57900 433629 57901
rect 433563 57836 433564 57900
rect 433628 57836 433629 57900
rect 433563 57835 433629 57836
rect 433379 57492 433445 57493
rect 433379 57428 433380 57492
rect 433444 57428 433445 57492
rect 433379 57427 433445 57428
rect 427675 57220 427741 57221
rect 427675 57156 427676 57220
rect 427740 57156 427741 57220
rect 427675 57155 427741 57156
rect 430987 57220 431053 57221
rect 430987 57156 430988 57220
rect 431052 57156 431053 57220
rect 430987 57155 431053 57156
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 434670 57901 434730 59470
rect 434667 57900 434733 57901
rect 434667 57836 434668 57900
rect 434732 57836 434733 57900
rect 434667 57835 434733 57836
rect 435774 57493 435834 59470
rect 435958 59470 436100 59530
rect 436878 59470 437052 59530
rect 438080 59530 438140 60106
rect 438488 59530 438548 60106
rect 439168 59530 439228 60106
rect 440936 59530 440996 60106
rect 443520 59530 443580 60106
rect 445968 59530 446028 60106
rect 438080 59470 438410 59530
rect 438488 59470 438594 59530
rect 435958 57901 436018 59470
rect 436878 57901 436938 59470
rect 435955 57900 436021 57901
rect 435955 57836 435956 57900
rect 436020 57836 436021 57900
rect 435955 57835 436021 57836
rect 436875 57900 436941 57901
rect 436875 57836 436876 57900
rect 436940 57836 436941 57900
rect 436875 57835 436941 57836
rect 435771 57492 435837 57493
rect 435771 57428 435772 57492
rect 435836 57428 435837 57492
rect 435771 57427 435837 57428
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 438350 57493 438410 59470
rect 438534 57901 438594 59470
rect 439086 59470 439228 59530
rect 440926 59470 440996 59530
rect 443502 59470 443580 59530
rect 445894 59470 446028 59530
rect 448280 59530 448340 60106
rect 451000 59530 451060 60106
rect 453448 59530 453508 60106
rect 455896 59530 455956 60106
rect 458480 59530 458540 60106
rect 448280 59470 448346 59530
rect 451000 59470 451106 59530
rect 438531 57900 438597 57901
rect 438531 57836 438532 57900
rect 438596 57836 438597 57900
rect 438531 57835 438597 57836
rect 438347 57492 438413 57493
rect 438347 57428 438348 57492
rect 438412 57428 438413 57492
rect 438347 57427 438413 57428
rect 439086 56269 439146 59470
rect 440926 57221 440986 59470
rect 440923 57220 440989 57221
rect 440923 57156 440924 57220
rect 440988 57156 440989 57220
rect 440923 57155 440989 57156
rect 439083 56268 439149 56269
rect 439083 56204 439084 56268
rect 439148 56204 439149 56268
rect 439083 56203 439149 56204
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 443502 57765 443562 59470
rect 443499 57764 443565 57765
rect 443499 57700 443500 57764
rect 443564 57700 443565 57764
rect 443499 57699 443565 57700
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 445894 57901 445954 59470
rect 445891 57900 445957 57901
rect 445891 57836 445892 57900
rect 445956 57836 445957 57900
rect 445891 57835 445957 57836
rect 448286 57357 448346 59470
rect 448283 57356 448349 57357
rect 448283 57292 448284 57356
rect 448348 57292 448349 57356
rect 448283 57291 448349 57292
rect 451046 56677 451106 59470
rect 453438 59470 453508 59530
rect 455830 59470 455956 59530
rect 458406 59470 458540 59530
rect 460928 59530 460988 60106
rect 463512 59530 463572 60106
rect 465960 59530 466020 60106
rect 468544 59530 468604 60106
rect 470992 59530 471052 60106
rect 460928 59470 461042 59530
rect 463512 59470 463618 59530
rect 453438 58853 453498 59470
rect 453435 58852 453501 58853
rect 453435 58788 453436 58852
rect 453500 58788 453501 58852
rect 453435 58787 453501 58788
rect 455830 58173 455890 59470
rect 458406 58581 458466 59470
rect 458403 58580 458469 58581
rect 458403 58516 458404 58580
rect 458468 58516 458469 58580
rect 458403 58515 458469 58516
rect 455827 58172 455893 58173
rect 455827 58108 455828 58172
rect 455892 58108 455893 58172
rect 455827 58107 455893 58108
rect 451794 57454 452414 58000
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451043 56676 451109 56677
rect 451043 56612 451044 56676
rect 451108 56612 451109 56676
rect 451043 56611 451109 56612
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 460982 57901 461042 59470
rect 463558 58717 463618 59470
rect 465950 59470 466020 59530
rect 468526 59470 468604 59530
rect 470918 59470 471052 59530
rect 473440 59530 473500 60106
rect 475888 59530 475948 60106
rect 478472 59530 478532 60106
rect 480920 59530 480980 60106
rect 473440 59470 473554 59530
rect 463555 58716 463621 58717
rect 463555 58652 463556 58716
rect 463620 58652 463621 58716
rect 463555 58651 463621 58652
rect 460979 57900 461045 57901
rect 460979 57836 460980 57900
rect 461044 57836 461045 57900
rect 460979 57835 461045 57836
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 465950 57901 466010 59470
rect 468526 58853 468586 59470
rect 468523 58852 468589 58853
rect 468523 58788 468524 58852
rect 468588 58788 468589 58852
rect 468523 58787 468589 58788
rect 465947 57900 466013 57901
rect 465947 57836 465948 57900
rect 466012 57836 466013 57900
rect 465947 57835 466013 57836
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 470918 57901 470978 59470
rect 473494 58989 473554 59470
rect 475886 59470 475948 59530
rect 478462 59470 478532 59530
rect 480854 59470 480980 59530
rect 483368 59530 483428 60106
rect 485952 59530 486012 60106
rect 503224 59530 503284 60106
rect 483368 59470 483490 59530
rect 485952 59470 486066 59530
rect 475886 58989 475946 59470
rect 473491 58988 473557 58989
rect 473491 58924 473492 58988
rect 473556 58924 473557 58988
rect 473491 58923 473557 58924
rect 475883 58988 475949 58989
rect 475883 58924 475884 58988
rect 475948 58924 475949 58988
rect 475883 58923 475949 58924
rect 470915 57900 470981 57901
rect 470915 57836 470916 57900
rect 470980 57836 470981 57900
rect 470915 57835 470981 57836
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 478462 57901 478522 59470
rect 480854 59261 480914 59470
rect 480851 59260 480917 59261
rect 480851 59196 480852 59260
rect 480916 59196 480917 59260
rect 480851 59195 480917 59196
rect 483430 59125 483490 59470
rect 483427 59124 483493 59125
rect 483427 59060 483428 59124
rect 483492 59060 483493 59124
rect 483427 59059 483493 59060
rect 478459 57900 478525 57901
rect 478459 57836 478460 57900
rect 478524 57836 478525 57900
rect 478459 57835 478525 57836
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 486006 57901 486066 59470
rect 503118 59470 503284 59530
rect 503360 59530 503420 60106
rect 503360 59470 503546 59530
rect 486003 57900 486069 57901
rect 486003 57836 486004 57900
rect 486068 57836 486069 57900
rect 486003 57835 486069 57836
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 503118 57901 503178 59470
rect 503486 57901 503546 59470
rect 503115 57900 503181 57901
rect 503115 57836 503116 57900
rect 503180 57836 503181 57900
rect 503115 57835 503181 57836
rect 503483 57900 503549 57901
rect 503483 57836 503484 57900
rect 503548 57836 503549 57900
rect 503483 57835 503549 57836
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 79610 597218 79846 597454
rect 79610 596898 79846 597134
rect 110330 597218 110566 597454
rect 110330 596898 110566 597134
rect 64250 579218 64486 579454
rect 64250 578898 64486 579134
rect 94970 579218 95206 579454
rect 94970 578898 95206 579134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 551598 63502 551834
rect 63586 551598 63822 551834
rect 63266 551278 63502 551514
rect 63586 551278 63822 551514
rect 66986 555318 67222 555554
rect 67306 555318 67542 555554
rect 66986 554998 67222 555234
rect 67306 554998 67542 555234
rect 73826 560278 74062 560514
rect 74146 560278 74382 560514
rect 73826 559958 74062 560194
rect 74146 559958 74382 560194
rect 77546 563998 77782 564234
rect 77866 563998 78102 564234
rect 77546 563678 77782 563914
rect 77866 563678 78102 563914
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 551598 99502 551834
rect 99586 551598 99822 551834
rect 99266 551278 99502 551514
rect 99586 551278 99822 551514
rect 102986 555318 103222 555554
rect 103306 555318 103542 555554
rect 102986 554998 103222 555234
rect 103306 554998 103542 555234
rect 109826 560278 110062 560514
rect 110146 560278 110382 560514
rect 109826 559958 110062 560194
rect 110146 559958 110382 560194
rect 113546 563998 113782 564234
rect 113866 563998 114102 564234
rect 113546 563678 113782 563914
rect 113866 563678 114102 563914
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 551598 135502 551834
rect 135586 551598 135822 551834
rect 135266 551278 135502 551514
rect 135586 551278 135822 551514
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 555318 139222 555554
rect 139306 555318 139542 555554
rect 138986 554998 139222 555234
rect 139306 554998 139542 555234
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 154250 615218 154486 615454
rect 154250 614898 154486 615134
rect 184970 615218 185206 615454
rect 184970 614898 185206 615134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 169610 597218 169846 597454
rect 169610 596898 169846 597134
rect 200330 597218 200566 597454
rect 200330 596898 200566 597134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 154250 579218 154486 579454
rect 154250 578898 154486 579134
rect 184970 579218 185206 579454
rect 184970 578898 185206 579134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 145826 560278 146062 560514
rect 146146 560278 146382 560514
rect 145826 559958 146062 560194
rect 146146 559958 146382 560194
rect 149546 563998 149782 564234
rect 149866 563998 150102 564234
rect 149546 563678 149782 563914
rect 149866 563678 150102 563914
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 551598 171502 551834
rect 171586 551598 171822 551834
rect 171266 551278 171502 551514
rect 171586 551278 171822 551514
rect 174986 555318 175222 555554
rect 175306 555318 175542 555554
rect 174986 554998 175222 555234
rect 175306 554998 175542 555234
rect 181826 560278 182062 560514
rect 182146 560278 182382 560514
rect 181826 559958 182062 560194
rect 182146 559958 182382 560194
rect 185546 563998 185782 564234
rect 185866 563998 186102 564234
rect 185546 563678 185782 563914
rect 185866 563678 186102 563914
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 551598 207502 551834
rect 207586 551598 207822 551834
rect 207266 551278 207502 551514
rect 207586 551278 207822 551514
rect 210986 555318 211222 555554
rect 211306 555318 211542 555554
rect 210986 554998 211222 555234
rect 211306 554998 211542 555234
rect 217826 560278 218062 560514
rect 218146 560278 218382 560514
rect 217826 559958 218062 560194
rect 218146 559958 218382 560194
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 563998 221782 564234
rect 221866 563998 222102 564234
rect 221546 563678 221782 563914
rect 221866 563678 222102 563914
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 244250 615218 244486 615454
rect 244250 614898 244486 615134
rect 274970 615218 275206 615454
rect 274970 614898 275206 615134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 259610 597218 259846 597454
rect 259610 596898 259846 597134
rect 290330 597218 290566 597454
rect 290330 596898 290566 597134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 244250 579218 244486 579454
rect 244250 578898 244486 579134
rect 274970 579218 275206 579454
rect 274970 578898 275206 579134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 551598 243502 551834
rect 243586 551598 243822 551834
rect 243266 551278 243502 551514
rect 243586 551278 243822 551514
rect 246986 555318 247222 555554
rect 247306 555318 247542 555554
rect 246986 554998 247222 555234
rect 247306 554998 247542 555234
rect 253826 560278 254062 560514
rect 254146 560278 254382 560514
rect 253826 559958 254062 560194
rect 254146 559958 254382 560194
rect 257546 563998 257782 564234
rect 257866 563998 258102 564234
rect 257546 563678 257782 563914
rect 257866 563678 258102 563914
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 551598 279502 551834
rect 279586 551598 279822 551834
rect 279266 551278 279502 551514
rect 279586 551278 279822 551514
rect 282986 555318 283222 555554
rect 283306 555318 283542 555554
rect 282986 554998 283222 555234
rect 283306 554998 283542 555234
rect 289826 560278 290062 560514
rect 290146 560278 290382 560514
rect 289826 559958 290062 560194
rect 290146 559958 290382 560194
rect 293546 563998 293782 564234
rect 293866 563998 294102 564234
rect 293546 563678 293782 563914
rect 293866 563678 294102 563914
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 64250 543218 64486 543454
rect 64250 542898 64486 543134
rect 94970 543218 95206 543454
rect 94970 542898 95206 543134
rect 125690 543218 125926 543454
rect 125690 542898 125926 543134
rect 156410 543218 156646 543454
rect 156410 542898 156646 543134
rect 187130 543218 187366 543454
rect 187130 542898 187366 543134
rect 217850 543218 218086 543454
rect 217850 542898 218086 543134
rect 248570 543218 248806 543454
rect 248570 542898 248806 543134
rect 279290 543218 279526 543454
rect 279290 542898 279526 543134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 79610 525218 79846 525454
rect 79610 524898 79846 525134
rect 110330 525218 110566 525454
rect 110330 524898 110566 525134
rect 141050 525218 141286 525454
rect 141050 524898 141286 525134
rect 171770 525218 172006 525454
rect 171770 524898 172006 525134
rect 202490 525218 202726 525454
rect 202490 524898 202726 525134
rect 233210 525218 233446 525454
rect 233210 524898 233446 525134
rect 263930 525218 264166 525454
rect 263930 524898 264166 525134
rect 294650 525218 294886 525454
rect 294650 524898 294886 525134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 475878 59782 476114
rect 59866 475878 60102 476114
rect 59546 475558 59782 475794
rect 59866 475558 60102 475794
rect 63266 477718 63502 477954
rect 63586 477718 63822 477954
rect 63266 477398 63502 477634
rect 63586 477398 63822 477634
rect 66986 481438 67222 481674
rect 67306 481438 67542 481674
rect 66986 481118 67222 481354
rect 67306 481118 67542 481354
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 472158 92062 472394
rect 92146 472158 92382 472394
rect 91826 471838 92062 472074
rect 92146 471838 92382 472074
rect 95546 475878 95782 476114
rect 95866 475878 96102 476114
rect 95546 475558 95782 475794
rect 95866 475558 96102 475794
rect 99266 477718 99502 477954
rect 99586 477718 99822 477954
rect 99266 477398 99502 477634
rect 99586 477398 99822 477634
rect 102986 481438 103222 481674
rect 103306 481438 103542 481674
rect 102986 481118 103222 481354
rect 103306 481118 103542 481354
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 472158 128062 472394
rect 128146 472158 128382 472394
rect 127826 471838 128062 472074
rect 128146 471838 128382 472074
rect 131546 475878 131782 476114
rect 131866 475878 132102 476114
rect 131546 475558 131782 475794
rect 131866 475558 132102 475794
rect 135266 477718 135502 477954
rect 135586 477718 135822 477954
rect 135266 477398 135502 477634
rect 135586 477398 135822 477634
rect 138986 481438 139222 481674
rect 139306 481438 139542 481674
rect 138986 481118 139222 481354
rect 139306 481118 139542 481354
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 472158 164062 472394
rect 164146 472158 164382 472394
rect 163826 471838 164062 472074
rect 164146 471838 164382 472074
rect 167546 475878 167782 476114
rect 167866 475878 168102 476114
rect 167546 475558 167782 475794
rect 167866 475558 168102 475794
rect 171266 477718 171502 477954
rect 171586 477718 171822 477954
rect 171266 477398 171502 477634
rect 171586 477398 171822 477634
rect 174986 481438 175222 481674
rect 175306 481438 175542 481674
rect 174986 481118 175222 481354
rect 175306 481118 175542 481354
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 61008 399218 61244 399454
rect 61008 398898 61244 399134
rect 195376 399218 195612 399454
rect 195376 398898 195612 399134
rect 59546 367878 59782 368114
rect 59866 367878 60102 368114
rect 59546 367558 59782 367794
rect 59866 367558 60102 367794
rect 63266 369718 63502 369954
rect 63586 369718 63822 369954
rect 63266 369398 63502 369634
rect 63586 369398 63822 369634
rect 66986 373438 67222 373674
rect 67306 373438 67542 373674
rect 66986 373118 67222 373354
rect 67306 373118 67542 373354
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 91826 364158 92062 364394
rect 92146 364158 92382 364394
rect 91826 363838 92062 364074
rect 92146 363838 92382 364074
rect 95546 367878 95782 368114
rect 95866 367878 96102 368114
rect 95546 367558 95782 367794
rect 95866 367558 96102 367794
rect 99266 369718 99502 369954
rect 99586 369718 99822 369954
rect 99266 369398 99502 369634
rect 99586 369398 99822 369634
rect 102986 373438 103222 373674
rect 103306 373438 103542 373674
rect 102986 373118 103222 373354
rect 103306 373118 103542 373354
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 364158 128062 364394
rect 128146 364158 128382 364394
rect 127826 363838 128062 364074
rect 128146 363838 128382 364074
rect 131546 367878 131782 368114
rect 131866 367878 132102 368114
rect 131546 367558 131782 367794
rect 131866 367558 132102 367794
rect 135266 369718 135502 369954
rect 135586 369718 135822 369954
rect 135266 369398 135502 369634
rect 135586 369398 135822 369634
rect 138986 373438 139222 373674
rect 139306 373438 139542 373674
rect 138986 373118 139222 373354
rect 139306 373118 139542 373354
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 163826 364158 164062 364394
rect 164146 364158 164382 364394
rect 163826 363838 164062 364074
rect 164146 363838 164382 364074
rect 167546 367878 167782 368114
rect 167866 367878 168102 368114
rect 167546 367558 167782 367794
rect 167866 367558 168102 367794
rect 171266 369718 171502 369954
rect 171586 369718 171822 369954
rect 171266 369398 171502 369634
rect 171586 369398 171822 369634
rect 174986 373438 175222 373674
rect 175306 373438 175542 373674
rect 174986 373118 175222 373354
rect 175306 373118 175542 373354
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 60328 345218 60564 345454
rect 60328 344898 60564 345134
rect 196056 345218 196292 345454
rect 196056 344898 196292 345134
rect 61008 327218 61244 327454
rect 61008 326898 61244 327134
rect 195376 327218 195612 327454
rect 195376 326898 195612 327134
rect 60328 309218 60564 309454
rect 60328 308898 60564 309134
rect 196056 309218 196292 309454
rect 196056 308898 196292 309134
rect 61008 291218 61244 291454
rect 61008 290898 61244 291134
rect 195376 291218 195612 291454
rect 195376 290898 195612 291134
rect 59546 259878 59782 260114
rect 59866 259878 60102 260114
rect 59546 259558 59782 259794
rect 59866 259558 60102 259794
rect 63266 261718 63502 261954
rect 63586 261718 63822 261954
rect 63266 261398 63502 261634
rect 63586 261398 63822 261634
rect 66986 265438 67222 265674
rect 67306 265438 67542 265674
rect 66986 265118 67222 265354
rect 67306 265118 67542 265354
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 91826 256158 92062 256394
rect 92146 256158 92382 256394
rect 91826 255838 92062 256074
rect 92146 255838 92382 256074
rect 95546 259878 95782 260114
rect 95866 259878 96102 260114
rect 95546 259558 95782 259794
rect 95866 259558 96102 259794
rect 99266 261718 99502 261954
rect 99586 261718 99822 261954
rect 99266 261398 99502 261634
rect 99586 261398 99822 261634
rect 102986 265438 103222 265674
rect 103306 265438 103542 265674
rect 102986 265118 103222 265354
rect 103306 265118 103542 265354
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 127826 256158 128062 256394
rect 128146 256158 128382 256394
rect 127826 255838 128062 256074
rect 128146 255838 128382 256074
rect 131546 259878 131782 260114
rect 131866 259878 132102 260114
rect 131546 259558 131782 259794
rect 131866 259558 132102 259794
rect 135266 261718 135502 261954
rect 135586 261718 135822 261954
rect 135266 261398 135502 261634
rect 135586 261398 135822 261634
rect 138986 265438 139222 265674
rect 139306 265438 139542 265674
rect 138986 265118 139222 265354
rect 139306 265118 139542 265354
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 256158 164062 256394
rect 164146 256158 164382 256394
rect 163826 255838 164062 256074
rect 164146 255838 164382 256074
rect 167546 259878 167782 260114
rect 167866 259878 168102 260114
rect 167546 259558 167782 259794
rect 167866 259558 168102 259794
rect 171266 261718 171502 261954
rect 171586 261718 171822 261954
rect 171266 261398 171502 261634
rect 171586 261398 171822 261634
rect 174986 265438 175222 265674
rect 175306 265438 175542 265674
rect 174986 265118 175222 265354
rect 175306 265118 175542 265354
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 60328 237218 60564 237454
rect 60328 236898 60564 237134
rect 196056 237218 196292 237454
rect 196056 236898 196292 237134
rect 61008 219218 61244 219454
rect 61008 218898 61244 219134
rect 195376 219218 195612 219454
rect 195376 218898 195612 219134
rect 60328 201218 60564 201454
rect 60328 200898 60564 201134
rect 196056 201218 196292 201454
rect 196056 200898 196292 201134
rect 61008 183218 61244 183454
rect 61008 182898 61244 183134
rect 195376 183218 195612 183454
rect 195376 182898 195612 183134
rect 59546 151878 59782 152114
rect 59866 151878 60102 152114
rect 59546 151558 59782 151794
rect 59866 151558 60102 151794
rect 63266 155598 63502 155834
rect 63586 155598 63822 155834
rect 63266 155278 63502 155514
rect 63586 155278 63822 155514
rect 66986 157438 67222 157674
rect 67306 157438 67542 157674
rect 66986 157118 67222 157354
rect 67306 157118 67542 157354
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 148158 92062 148394
rect 92146 148158 92382 148394
rect 91826 147838 92062 148074
rect 92146 147838 92382 148074
rect 95546 151878 95782 152114
rect 95866 151878 96102 152114
rect 95546 151558 95782 151794
rect 95866 151558 96102 151794
rect 99266 155598 99502 155834
rect 99586 155598 99822 155834
rect 99266 155278 99502 155514
rect 99586 155278 99822 155514
rect 102986 157438 103222 157674
rect 103306 157438 103542 157674
rect 102986 157118 103222 157354
rect 103306 157118 103542 157354
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 127826 148158 128062 148394
rect 128146 148158 128382 148394
rect 127826 147838 128062 148074
rect 128146 147838 128382 148074
rect 131546 151878 131782 152114
rect 131866 151878 132102 152114
rect 131546 151558 131782 151794
rect 131866 151558 132102 151794
rect 135266 155598 135502 155834
rect 135586 155598 135822 155834
rect 135266 155278 135502 155514
rect 135586 155278 135822 155514
rect 138986 157438 139222 157674
rect 139306 157438 139542 157674
rect 138986 157118 139222 157354
rect 139306 157118 139542 157354
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 163826 148158 164062 148394
rect 164146 148158 164382 148394
rect 163826 147838 164062 148074
rect 164146 147838 164382 148074
rect 167546 151878 167782 152114
rect 167866 151878 168102 152114
rect 167546 151558 167782 151794
rect 167866 151558 168102 151794
rect 171266 155598 171502 155834
rect 171586 155598 171822 155834
rect 171266 155278 171502 155514
rect 171586 155278 171822 155514
rect 174986 157438 175222 157674
rect 175306 157438 175542 157674
rect 174986 157118 175222 157354
rect 175306 157118 175542 157354
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 60328 129218 60564 129454
rect 60328 128898 60564 129134
rect 196056 129218 196292 129454
rect 196056 128898 196292 129134
rect 61008 111218 61244 111454
rect 61008 110898 61244 111134
rect 195376 111218 195612 111454
rect 195376 110898 195612 111134
rect 60328 93218 60564 93454
rect 60328 92898 60564 93134
rect 196056 93218 196292 93454
rect 196056 92898 196292 93134
rect 61008 75218 61244 75454
rect 61008 74898 61244 75134
rect 195376 75218 195612 75454
rect 195376 74898 195612 75134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 199826 472158 200062 472394
rect 200146 472158 200382 472394
rect 199826 471838 200062 472074
rect 200146 471838 200382 472074
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 364158 200062 364394
rect 200146 364158 200382 364394
rect 199826 363838 200062 364074
rect 200146 363838 200382 364074
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 256158 200062 256394
rect 200146 256158 200382 256394
rect 199826 255838 200062 256074
rect 200146 255838 200382 256074
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 148158 200062 148394
rect 200146 148158 200382 148394
rect 199826 147838 200062 148074
rect 200146 147838 200382 148074
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 203546 475878 203782 476114
rect 203866 475878 204102 476114
rect 203546 475558 203782 475794
rect 203866 475558 204102 475794
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 367878 203782 368114
rect 203866 367878 204102 368114
rect 203546 367558 203782 367794
rect 203866 367558 204102 367794
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 259878 203782 260114
rect 203866 259878 204102 260114
rect 203546 259558 203782 259794
rect 203866 259558 204102 259794
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 151878 203782 152114
rect 203866 151878 204102 152114
rect 203546 151558 203782 151794
rect 203866 151558 204102 151794
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 207266 477718 207502 477954
rect 207586 477718 207822 477954
rect 207266 477398 207502 477634
rect 207586 477398 207822 477634
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 369718 207502 369954
rect 207586 369718 207822 369954
rect 207266 369398 207502 369634
rect 207586 369398 207822 369634
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 261718 207502 261954
rect 207586 261718 207822 261954
rect 207266 261398 207502 261634
rect 207586 261398 207822 261634
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 210986 481438 211222 481674
rect 211306 481438 211542 481674
rect 210986 481118 211222 481354
rect 211306 481118 211542 481354
rect 207266 155598 207502 155834
rect 207586 155598 207822 155834
rect 207266 155278 207502 155514
rect 207586 155278 207822 155514
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 373438 211222 373674
rect 211306 373438 211542 373674
rect 210986 373118 211222 373354
rect 211306 373118 211542 373354
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 265438 211222 265674
rect 211306 265438 211542 265674
rect 210986 265118 211222 265354
rect 211306 265118 211542 265354
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 157438 211222 157674
rect 211306 157438 211542 157674
rect 210986 157118 211222 157354
rect 211306 157118 211542 157354
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 472158 236062 472394
rect 236146 472158 236382 472394
rect 235826 471838 236062 472074
rect 236146 471838 236382 472074
rect 239546 475878 239782 476114
rect 239866 475878 240102 476114
rect 239546 475558 239782 475794
rect 239866 475558 240102 475794
rect 243266 477718 243502 477954
rect 243586 477718 243822 477954
rect 243266 477398 243502 477634
rect 243586 477398 243822 477634
rect 246986 481438 247222 481674
rect 247306 481438 247542 481674
rect 246986 481118 247222 481354
rect 247306 481118 247542 481354
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 472158 272062 472394
rect 272146 472158 272382 472394
rect 271826 471838 272062 472074
rect 272146 471838 272382 472074
rect 275546 475878 275782 476114
rect 275866 475878 276102 476114
rect 275546 475558 275782 475794
rect 275866 475558 276102 475794
rect 279266 477718 279502 477954
rect 279586 477718 279822 477954
rect 279266 477398 279502 477634
rect 279586 477398 279822 477634
rect 282986 481438 283222 481674
rect 283306 481438 283542 481674
rect 282986 481118 283222 481354
rect 283306 481118 283542 481354
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 329250 615218 329486 615454
rect 329250 614898 329486 615134
rect 359970 615218 360206 615454
rect 359970 614898 360206 615134
rect 390690 615218 390926 615454
rect 390690 614898 390926 615134
rect 421410 615218 421646 615454
rect 421410 614898 421646 615134
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 344610 597218 344846 597454
rect 344610 596898 344846 597134
rect 375330 597218 375566 597454
rect 375330 596898 375566 597134
rect 406050 597218 406286 597454
rect 406050 596898 406286 597134
rect 329250 579218 329486 579454
rect 329250 578898 329486 579134
rect 359970 579218 360206 579454
rect 359970 578898 360206 579134
rect 390690 579218 390926 579454
rect 390690 578898 390926 579134
rect 421410 579218 421646 579454
rect 421410 578898 421646 579134
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 344610 561218 344846 561454
rect 344610 560898 344846 561134
rect 375330 561218 375566 561454
rect 375330 560898 375566 561134
rect 406050 561218 406286 561454
rect 406050 560898 406286 561134
rect 329250 543218 329486 543454
rect 329250 542898 329486 543134
rect 359970 543218 360206 543454
rect 359970 542898 360206 543134
rect 390690 543218 390926 543454
rect 390690 542898 390926 543134
rect 421410 543218 421646 543454
rect 421410 542898 421646 543134
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 344610 525218 344846 525454
rect 344610 524898 344846 525134
rect 375330 525218 375566 525454
rect 375330 524898 375566 525134
rect 406050 525218 406286 525454
rect 406050 524898 406286 525134
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221008 399218 221244 399454
rect 221008 398898 221244 399134
rect 355376 399218 355612 399454
rect 355376 398898 355612 399134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 364158 236062 364394
rect 236146 364158 236382 364394
rect 235826 363838 236062 364074
rect 236146 363838 236382 364074
rect 239546 367878 239782 368114
rect 239866 367878 240102 368114
rect 239546 367558 239782 367794
rect 239866 367558 240102 367794
rect 243266 369718 243502 369954
rect 243586 369718 243822 369954
rect 243266 369398 243502 369634
rect 243586 369398 243822 369634
rect 246986 373438 247222 373674
rect 247306 373438 247542 373674
rect 246986 373118 247222 373354
rect 247306 373118 247542 373354
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 364158 272062 364394
rect 272146 364158 272382 364394
rect 271826 363838 272062 364074
rect 272146 363838 272382 364074
rect 275546 367878 275782 368114
rect 275866 367878 276102 368114
rect 275546 367558 275782 367794
rect 275866 367558 276102 367794
rect 279266 369718 279502 369954
rect 279586 369718 279822 369954
rect 279266 369398 279502 369634
rect 279586 369398 279822 369634
rect 282986 373438 283222 373674
rect 283306 373438 283542 373674
rect 282986 373118 283222 373354
rect 283306 373118 283542 373354
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 364158 308062 364394
rect 308146 364158 308382 364394
rect 307826 363838 308062 364074
rect 308146 363838 308382 364074
rect 311546 367878 311782 368114
rect 311866 367878 312102 368114
rect 311546 367558 311782 367794
rect 311866 367558 312102 367794
rect 315266 369718 315502 369954
rect 315586 369718 315822 369954
rect 315266 369398 315502 369634
rect 315586 369398 315822 369634
rect 318986 373438 319222 373674
rect 319306 373438 319542 373674
rect 318986 373118 319222 373354
rect 319306 373118 319542 373354
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 343826 364158 344062 364394
rect 344146 364158 344382 364394
rect 343826 363838 344062 364074
rect 344146 363838 344382 364074
rect 347546 367878 347782 368114
rect 347866 367878 348102 368114
rect 347546 367558 347782 367794
rect 347866 367558 348102 367794
rect 351266 369718 351502 369954
rect 351586 369718 351822 369954
rect 351266 369398 351502 369634
rect 351586 369398 351822 369634
rect 354986 373438 355222 373674
rect 355306 373438 355542 373674
rect 354986 373118 355222 373354
rect 355306 373118 355542 373354
rect 220328 345218 220564 345454
rect 220328 344898 220564 345134
rect 356056 345218 356292 345454
rect 356056 344898 356292 345134
rect 221008 327218 221244 327454
rect 221008 326898 221244 327134
rect 355376 327218 355612 327454
rect 355376 326898 355612 327134
rect 220328 309218 220564 309454
rect 220328 308898 220564 309134
rect 356056 309218 356292 309454
rect 356056 308898 356292 309134
rect 221008 291218 221244 291454
rect 221008 290898 221244 291134
rect 355376 291218 355612 291454
rect 355376 290898 355612 291134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 235826 256158 236062 256394
rect 236146 256158 236382 256394
rect 235826 255838 236062 256074
rect 236146 255838 236382 256074
rect 239546 259878 239782 260114
rect 239866 259878 240102 260114
rect 239546 259558 239782 259794
rect 239866 259558 240102 259794
rect 243266 261718 243502 261954
rect 243586 261718 243822 261954
rect 243266 261398 243502 261634
rect 243586 261398 243822 261634
rect 246986 265438 247222 265674
rect 247306 265438 247542 265674
rect 246986 265118 247222 265354
rect 247306 265118 247542 265354
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 271826 256158 272062 256394
rect 272146 256158 272382 256394
rect 271826 255838 272062 256074
rect 272146 255838 272382 256074
rect 275546 259878 275782 260114
rect 275866 259878 276102 260114
rect 275546 259558 275782 259794
rect 275866 259558 276102 259794
rect 279266 261718 279502 261954
rect 279586 261718 279822 261954
rect 279266 261398 279502 261634
rect 279586 261398 279822 261634
rect 282986 265438 283222 265674
rect 283306 265438 283542 265674
rect 282986 265118 283222 265354
rect 283306 265118 283542 265354
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 307826 256158 308062 256394
rect 308146 256158 308382 256394
rect 307826 255838 308062 256074
rect 308146 255838 308382 256074
rect 311546 259878 311782 260114
rect 311866 259878 312102 260114
rect 311546 259558 311782 259794
rect 311866 259558 312102 259794
rect 315266 261718 315502 261954
rect 315586 261718 315822 261954
rect 315266 261398 315502 261634
rect 315586 261398 315822 261634
rect 318986 265438 319222 265674
rect 319306 265438 319542 265674
rect 318986 265118 319222 265354
rect 319306 265118 319542 265354
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 343826 256158 344062 256394
rect 344146 256158 344382 256394
rect 343826 255838 344062 256074
rect 344146 255838 344382 256074
rect 347546 259878 347782 260114
rect 347866 259878 348102 260114
rect 347546 259558 347782 259794
rect 347866 259558 348102 259794
rect 351266 261718 351502 261954
rect 351586 261718 351822 261954
rect 351266 261398 351502 261634
rect 351586 261398 351822 261634
rect 354986 265438 355222 265674
rect 355306 265438 355542 265674
rect 354986 265118 355222 265354
rect 355306 265118 355542 265354
rect 220328 237218 220564 237454
rect 220328 236898 220564 237134
rect 356056 237218 356292 237454
rect 356056 236898 356292 237134
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 201218 220564 201454
rect 220328 200898 220564 201134
rect 356056 201218 356292 201454
rect 356056 200898 356292 201134
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 235826 148158 236062 148394
rect 236146 148158 236382 148394
rect 235826 147838 236062 148074
rect 236146 147838 236382 148074
rect 239546 151878 239782 152114
rect 239866 151878 240102 152114
rect 239546 151558 239782 151794
rect 239866 151558 240102 151794
rect 243266 155598 243502 155834
rect 243586 155598 243822 155834
rect 243266 155278 243502 155514
rect 243586 155278 243822 155514
rect 246986 157438 247222 157674
rect 247306 157438 247542 157674
rect 246986 157118 247222 157354
rect 247306 157118 247542 157354
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 271826 148158 272062 148394
rect 272146 148158 272382 148394
rect 271826 147838 272062 148074
rect 272146 147838 272382 148074
rect 275546 151878 275782 152114
rect 275866 151878 276102 152114
rect 275546 151558 275782 151794
rect 275866 151558 276102 151794
rect 279266 155598 279502 155834
rect 279586 155598 279822 155834
rect 279266 155278 279502 155514
rect 279586 155278 279822 155514
rect 282986 157438 283222 157674
rect 283306 157438 283542 157674
rect 282986 157118 283222 157354
rect 283306 157118 283542 157354
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 307826 148158 308062 148394
rect 308146 148158 308382 148394
rect 307826 147838 308062 148074
rect 308146 147838 308382 148074
rect 311546 151878 311782 152114
rect 311866 151878 312102 152114
rect 311546 151558 311782 151794
rect 311866 151558 312102 151794
rect 315266 155598 315502 155834
rect 315586 155598 315822 155834
rect 315266 155278 315502 155514
rect 315586 155278 315822 155514
rect 318986 157438 319222 157674
rect 319306 157438 319542 157674
rect 318986 157118 319222 157354
rect 319306 157118 319542 157354
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 343826 148158 344062 148394
rect 344146 148158 344382 148394
rect 343826 147838 344062 148074
rect 344146 147838 344382 148074
rect 347546 151878 347782 152114
rect 347866 151878 348102 152114
rect 347546 151558 347782 151794
rect 347866 151558 348102 151794
rect 351266 155598 351502 155834
rect 351586 155598 351822 155834
rect 351266 155278 351502 155514
rect 351586 155278 351822 155514
rect 354986 157438 355222 157674
rect 355306 157438 355542 157674
rect 354986 157118 355222 157354
rect 355306 157118 355542 157354
rect 220328 129218 220564 129454
rect 220328 128898 220564 129134
rect 356056 129218 356292 129454
rect 356056 128898 356292 129134
rect 221008 111218 221244 111454
rect 221008 110898 221244 111134
rect 355376 111218 355612 111454
rect 355376 110898 355612 111134
rect 220328 93218 220564 93454
rect 220328 92898 220564 93134
rect 356056 93218 356292 93454
rect 356056 92898 356292 93134
rect 221008 75218 221244 75454
rect 221008 74898 221244 75134
rect 355376 75218 355612 75454
rect 355376 74898 355612 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 479610 597218 479846 597454
rect 479610 596898 479846 597134
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 380328 453218 380564 453454
rect 380328 452898 380564 453134
rect 516056 453218 516292 453454
rect 516056 452898 516292 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 381008 435218 381244 435454
rect 381008 434898 381244 435134
rect 515376 435218 515612 435454
rect 515376 434898 515612 435134
rect 380328 417218 380564 417454
rect 380328 416898 380564 417134
rect 516056 417218 516292 417454
rect 516056 416898 516292 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 381008 399218 381244 399454
rect 381008 398898 381244 399134
rect 515376 399218 515612 399454
rect 515376 398898 515612 399134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 379826 364158 380062 364394
rect 380146 364158 380382 364394
rect 379826 363838 380062 364074
rect 380146 363838 380382 364074
rect 383546 367878 383782 368114
rect 383866 367878 384102 368114
rect 383546 367558 383782 367794
rect 383866 367558 384102 367794
rect 387266 369718 387502 369954
rect 387586 369718 387822 369954
rect 387266 369398 387502 369634
rect 387586 369398 387822 369634
rect 390986 373438 391222 373674
rect 391306 373438 391542 373674
rect 390986 373118 391222 373354
rect 391306 373118 391542 373354
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 415826 364158 416062 364394
rect 416146 364158 416382 364394
rect 415826 363838 416062 364074
rect 416146 363838 416382 364074
rect 419546 367878 419782 368114
rect 419866 367878 420102 368114
rect 419546 367558 419782 367794
rect 419866 367558 420102 367794
rect 423266 369718 423502 369954
rect 423586 369718 423822 369954
rect 423266 369398 423502 369634
rect 423586 369398 423822 369634
rect 426986 373438 427222 373674
rect 427306 373438 427542 373674
rect 426986 373118 427222 373354
rect 427306 373118 427542 373354
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 451826 364158 452062 364394
rect 452146 364158 452382 364394
rect 451826 363838 452062 364074
rect 452146 363838 452382 364074
rect 455546 367878 455782 368114
rect 455866 367878 456102 368114
rect 455546 367558 455782 367794
rect 455866 367558 456102 367794
rect 459266 369718 459502 369954
rect 459586 369718 459822 369954
rect 459266 369398 459502 369634
rect 459586 369398 459822 369634
rect 462986 373438 463222 373674
rect 463306 373438 463542 373674
rect 462986 373118 463222 373354
rect 463306 373118 463542 373354
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 487826 364158 488062 364394
rect 488146 364158 488382 364394
rect 487826 363838 488062 364074
rect 488146 363838 488382 364074
rect 491546 367878 491782 368114
rect 491866 367878 492102 368114
rect 491546 367558 491782 367794
rect 491866 367558 492102 367794
rect 495266 369718 495502 369954
rect 495586 369718 495822 369954
rect 495266 369398 495502 369634
rect 495586 369398 495822 369634
rect 498986 373438 499222 373674
rect 499306 373438 499542 373674
rect 498986 373118 499222 373354
rect 499306 373118 499542 373354
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 380328 345218 380564 345454
rect 380328 344898 380564 345134
rect 516056 345218 516292 345454
rect 516056 344898 516292 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 381008 327218 381244 327454
rect 381008 326898 381244 327134
rect 515376 327218 515612 327454
rect 515376 326898 515612 327134
rect 380328 309218 380564 309454
rect 380328 308898 380564 309134
rect 516056 309218 516292 309454
rect 516056 308898 516292 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 381008 291218 381244 291454
rect 381008 290898 381244 291134
rect 515376 291218 515612 291454
rect 515376 290898 515612 291134
rect 379826 256158 380062 256394
rect 380146 256158 380382 256394
rect 379826 255838 380062 256074
rect 380146 255838 380382 256074
rect 383546 259878 383782 260114
rect 383866 259878 384102 260114
rect 383546 259558 383782 259794
rect 383866 259558 384102 259794
rect 387266 261718 387502 261954
rect 387586 261718 387822 261954
rect 387266 261398 387502 261634
rect 387586 261398 387822 261634
rect 390986 265438 391222 265674
rect 391306 265438 391542 265674
rect 390986 265118 391222 265354
rect 391306 265118 391542 265354
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 415826 256158 416062 256394
rect 416146 256158 416382 256394
rect 415826 255838 416062 256074
rect 416146 255838 416382 256074
rect 419546 259878 419782 260114
rect 419866 259878 420102 260114
rect 419546 259558 419782 259794
rect 419866 259558 420102 259794
rect 423266 261718 423502 261954
rect 423586 261718 423822 261954
rect 423266 261398 423502 261634
rect 423586 261398 423822 261634
rect 426986 265438 427222 265674
rect 427306 265438 427542 265674
rect 426986 265118 427222 265354
rect 427306 265118 427542 265354
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 451826 256158 452062 256394
rect 452146 256158 452382 256394
rect 451826 255838 452062 256074
rect 452146 255838 452382 256074
rect 455546 259878 455782 260114
rect 455866 259878 456102 260114
rect 455546 259558 455782 259794
rect 455866 259558 456102 259794
rect 459266 261718 459502 261954
rect 459586 261718 459822 261954
rect 459266 261398 459502 261634
rect 459586 261398 459822 261634
rect 462986 265438 463222 265674
rect 463306 265438 463542 265674
rect 462986 265118 463222 265354
rect 463306 265118 463542 265354
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 487826 256158 488062 256394
rect 488146 256158 488382 256394
rect 487826 255838 488062 256074
rect 488146 255838 488382 256074
rect 491546 259878 491782 260114
rect 491866 259878 492102 260114
rect 491546 259558 491782 259794
rect 491866 259558 492102 259794
rect 495266 261718 495502 261954
rect 495586 261718 495822 261954
rect 495266 261398 495502 261634
rect 495586 261398 495822 261634
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 498986 265438 499222 265674
rect 499306 265438 499542 265674
rect 498986 265118 499222 265354
rect 499306 265118 499542 265354
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 380328 237218 380564 237454
rect 380328 236898 380564 237134
rect 516056 237218 516292 237454
rect 516056 236898 516292 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 381008 219218 381244 219454
rect 381008 218898 381244 219134
rect 515376 219218 515612 219454
rect 515376 218898 515612 219134
rect 380328 201218 380564 201454
rect 380328 200898 380564 201134
rect 516056 201218 516292 201454
rect 516056 200898 516292 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 381008 183218 381244 183454
rect 381008 182898 381244 183134
rect 515376 183218 515612 183454
rect 515376 182898 515612 183134
rect 379826 148158 380062 148394
rect 380146 148158 380382 148394
rect 379826 147838 380062 148074
rect 380146 147838 380382 148074
rect 383546 151878 383782 152114
rect 383866 151878 384102 152114
rect 383546 151558 383782 151794
rect 383866 151558 384102 151794
rect 387266 155598 387502 155834
rect 387586 155598 387822 155834
rect 387266 155278 387502 155514
rect 387586 155278 387822 155514
rect 390986 157438 391222 157674
rect 391306 157438 391542 157674
rect 390986 157118 391222 157354
rect 391306 157118 391542 157354
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 415826 148158 416062 148394
rect 416146 148158 416382 148394
rect 415826 147838 416062 148074
rect 416146 147838 416382 148074
rect 419546 151878 419782 152114
rect 419866 151878 420102 152114
rect 419546 151558 419782 151794
rect 419866 151558 420102 151794
rect 423266 155598 423502 155834
rect 423586 155598 423822 155834
rect 423266 155278 423502 155514
rect 423586 155278 423822 155514
rect 426986 157438 427222 157674
rect 427306 157438 427542 157674
rect 426986 157118 427222 157354
rect 427306 157118 427542 157354
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 148158 452062 148394
rect 452146 148158 452382 148394
rect 451826 147838 452062 148074
rect 452146 147838 452382 148074
rect 455546 151878 455782 152114
rect 455866 151878 456102 152114
rect 455546 151558 455782 151794
rect 455866 151558 456102 151794
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 459266 155598 459502 155834
rect 459586 155598 459822 155834
rect 459266 155278 459502 155514
rect 459586 155278 459822 155514
rect 462986 157438 463222 157674
rect 463306 157438 463542 157674
rect 462986 157118 463222 157354
rect 463306 157118 463542 157354
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 148158 488062 148394
rect 488146 148158 488382 148394
rect 487826 147838 488062 148074
rect 488146 147838 488382 148074
rect 491546 151878 491782 152114
rect 491866 151878 492102 152114
rect 491546 151558 491782 151794
rect 491866 151558 492102 151794
rect 495266 155598 495502 155834
rect 495586 155598 495822 155834
rect 495266 155278 495502 155514
rect 495586 155278 495822 155514
rect 498986 157438 499222 157674
rect 499306 157438 499542 157674
rect 498986 157118 499222 157354
rect 499306 157118 499542 157354
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 380328 129218 380564 129454
rect 380328 128898 380564 129134
rect 516056 129218 516292 129454
rect 516056 128898 516292 129134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 381008 111218 381244 111454
rect 381008 110898 381244 111134
rect 515376 111218 515612 111454
rect 515376 110898 515612 111134
rect 380328 93218 380564 93454
rect 380328 92898 380564 93134
rect 516056 93218 516292 93454
rect 516056 92898 516292 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 381008 75218 381244 75454
rect 381008 74898 381244 75134
rect 515376 75218 515612 75454
rect 515376 74898 515612 75134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 154250 615454
rect 154486 615218 184970 615454
rect 185206 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 244250 615454
rect 244486 615218 274970 615454
rect 275206 615218 329250 615454
rect 329486 615218 359970 615454
rect 360206 615218 390690 615454
rect 390926 615218 421410 615454
rect 421646 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 154250 615134
rect 154486 614898 184970 615134
rect 185206 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 244250 615134
rect 244486 614898 274970 615134
rect 275206 614898 329250 615134
rect 329486 614898 359970 615134
rect 360206 614898 390690 615134
rect 390926 614898 421410 615134
rect 421646 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 79610 597454
rect 79846 597218 110330 597454
rect 110566 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 169610 597454
rect 169846 597218 200330 597454
rect 200566 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 259610 597454
rect 259846 597218 290330 597454
rect 290566 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 344610 597454
rect 344846 597218 375330 597454
rect 375566 597218 406050 597454
rect 406286 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 479610 597454
rect 479846 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 79610 597134
rect 79846 596898 110330 597134
rect 110566 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 169610 597134
rect 169846 596898 200330 597134
rect 200566 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 259610 597134
rect 259846 596898 290330 597134
rect 290566 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 344610 597134
rect 344846 596898 375330 597134
rect 375566 596898 406050 597134
rect 406286 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 479610 597134
rect 479846 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64250 579454
rect 64486 579218 94970 579454
rect 95206 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 154250 579454
rect 154486 579218 184970 579454
rect 185206 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 244250 579454
rect 244486 579218 274970 579454
rect 275206 579218 329250 579454
rect 329486 579218 359970 579454
rect 360206 579218 390690 579454
rect 390926 579218 421410 579454
rect 421646 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64250 579134
rect 64486 578898 94970 579134
rect 95206 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 154250 579134
rect 154486 578898 184970 579134
rect 185206 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 244250 579134
rect 244486 578898 274970 579134
rect 275206 578898 329250 579134
rect 329486 578898 359970 579134
rect 360206 578898 390690 579134
rect 390926 578898 421410 579134
rect 421646 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect 77514 564234 294134 564266
rect 77514 563998 77546 564234
rect 77782 563998 77866 564234
rect 78102 563998 113546 564234
rect 113782 563998 113866 564234
rect 114102 563998 149546 564234
rect 149782 563998 149866 564234
rect 150102 563998 185546 564234
rect 185782 563998 185866 564234
rect 186102 563998 221546 564234
rect 221782 563998 221866 564234
rect 222102 563998 257546 564234
rect 257782 563998 257866 564234
rect 258102 563998 293546 564234
rect 293782 563998 293866 564234
rect 294102 563998 294134 564234
rect 77514 563914 294134 563998
rect 77514 563678 77546 563914
rect 77782 563678 77866 563914
rect 78102 563678 113546 563914
rect 113782 563678 113866 563914
rect 114102 563678 149546 563914
rect 149782 563678 149866 563914
rect 150102 563678 185546 563914
rect 185782 563678 185866 563914
rect 186102 563678 221546 563914
rect 221782 563678 221866 563914
rect 222102 563678 257546 563914
rect 257782 563678 257866 563914
rect 258102 563678 293546 563914
rect 293782 563678 293866 563914
rect 294102 563678 294134 563914
rect 77514 563646 294134 563678
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 344610 561454
rect 344846 561218 375330 561454
rect 375566 561218 406050 561454
rect 406286 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 344610 561134
rect 344846 560898 375330 561134
rect 375566 560898 406050 561134
rect 406286 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect 73794 560514 290414 560546
rect 73794 560278 73826 560514
rect 74062 560278 74146 560514
rect 74382 560278 109826 560514
rect 110062 560278 110146 560514
rect 110382 560278 145826 560514
rect 146062 560278 146146 560514
rect 146382 560278 181826 560514
rect 182062 560278 182146 560514
rect 182382 560278 217826 560514
rect 218062 560278 218146 560514
rect 218382 560278 253826 560514
rect 254062 560278 254146 560514
rect 254382 560278 289826 560514
rect 290062 560278 290146 560514
rect 290382 560278 290414 560514
rect 73794 560194 290414 560278
rect 73794 559958 73826 560194
rect 74062 559958 74146 560194
rect 74382 559958 109826 560194
rect 110062 559958 110146 560194
rect 110382 559958 145826 560194
rect 146062 559958 146146 560194
rect 146382 559958 181826 560194
rect 182062 559958 182146 560194
rect 182382 559958 217826 560194
rect 218062 559958 218146 560194
rect 218382 559958 253826 560194
rect 254062 559958 254146 560194
rect 254382 559958 289826 560194
rect 290062 559958 290146 560194
rect 290382 559958 290414 560194
rect 73794 559926 290414 559958
rect 66954 555554 283574 555586
rect 66954 555318 66986 555554
rect 67222 555318 67306 555554
rect 67542 555318 102986 555554
rect 103222 555318 103306 555554
rect 103542 555318 138986 555554
rect 139222 555318 139306 555554
rect 139542 555318 174986 555554
rect 175222 555318 175306 555554
rect 175542 555318 210986 555554
rect 211222 555318 211306 555554
rect 211542 555318 246986 555554
rect 247222 555318 247306 555554
rect 247542 555318 282986 555554
rect 283222 555318 283306 555554
rect 283542 555318 283574 555554
rect 66954 555234 283574 555318
rect 66954 554998 66986 555234
rect 67222 554998 67306 555234
rect 67542 554998 102986 555234
rect 103222 554998 103306 555234
rect 103542 554998 138986 555234
rect 139222 554998 139306 555234
rect 139542 554998 174986 555234
rect 175222 554998 175306 555234
rect 175542 554998 210986 555234
rect 211222 554998 211306 555234
rect 211542 554998 246986 555234
rect 247222 554998 247306 555234
rect 247542 554998 282986 555234
rect 283222 554998 283306 555234
rect 283542 554998 283574 555234
rect 66954 554966 283574 554998
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect 63234 551834 279854 551866
rect 63234 551598 63266 551834
rect 63502 551598 63586 551834
rect 63822 551598 99266 551834
rect 99502 551598 99586 551834
rect 99822 551598 135266 551834
rect 135502 551598 135586 551834
rect 135822 551598 171266 551834
rect 171502 551598 171586 551834
rect 171822 551598 207266 551834
rect 207502 551598 207586 551834
rect 207822 551598 243266 551834
rect 243502 551598 243586 551834
rect 243822 551598 279266 551834
rect 279502 551598 279586 551834
rect 279822 551598 279854 551834
rect 63234 551514 279854 551598
rect 63234 551278 63266 551514
rect 63502 551278 63586 551514
rect 63822 551278 99266 551514
rect 99502 551278 99586 551514
rect 99822 551278 135266 551514
rect 135502 551278 135586 551514
rect 135822 551278 171266 551514
rect 171502 551278 171586 551514
rect 171822 551278 207266 551514
rect 207502 551278 207586 551514
rect 207822 551278 243266 551514
rect 243502 551278 243586 551514
rect 243822 551278 279266 551514
rect 279502 551278 279586 551514
rect 279822 551278 279854 551514
rect 63234 551246 279854 551278
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 64250 543454
rect 64486 543218 94970 543454
rect 95206 543218 125690 543454
rect 125926 543218 156410 543454
rect 156646 543218 187130 543454
rect 187366 543218 217850 543454
rect 218086 543218 248570 543454
rect 248806 543218 279290 543454
rect 279526 543218 329250 543454
rect 329486 543218 359970 543454
rect 360206 543218 390690 543454
rect 390926 543218 421410 543454
rect 421646 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 64250 543134
rect 64486 542898 94970 543134
rect 95206 542898 125690 543134
rect 125926 542898 156410 543134
rect 156646 542898 187130 543134
rect 187366 542898 217850 543134
rect 218086 542898 248570 543134
rect 248806 542898 279290 543134
rect 279526 542898 329250 543134
rect 329486 542898 359970 543134
rect 360206 542898 390690 543134
rect 390926 542898 421410 543134
rect 421646 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 79610 525454
rect 79846 525218 110330 525454
rect 110566 525218 141050 525454
rect 141286 525218 171770 525454
rect 172006 525218 202490 525454
rect 202726 525218 233210 525454
rect 233446 525218 263930 525454
rect 264166 525218 294650 525454
rect 294886 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 344610 525454
rect 344846 525218 375330 525454
rect 375566 525218 406050 525454
rect 406286 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 79610 525134
rect 79846 524898 110330 525134
rect 110566 524898 141050 525134
rect 141286 524898 171770 525134
rect 172006 524898 202490 525134
rect 202726 524898 233210 525134
rect 233446 524898 263930 525134
rect 264166 524898 294650 525134
rect 294886 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 344610 525134
rect 344846 524898 375330 525134
rect 375566 524898 406050 525134
rect 406286 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect 66954 481674 283574 481706
rect 66954 481438 66986 481674
rect 67222 481438 67306 481674
rect 67542 481438 102986 481674
rect 103222 481438 103306 481674
rect 103542 481438 138986 481674
rect 139222 481438 139306 481674
rect 139542 481438 174986 481674
rect 175222 481438 175306 481674
rect 175542 481438 210986 481674
rect 211222 481438 211306 481674
rect 211542 481438 246986 481674
rect 247222 481438 247306 481674
rect 247542 481438 282986 481674
rect 283222 481438 283306 481674
rect 283542 481438 283574 481674
rect 66954 481354 283574 481438
rect 66954 481118 66986 481354
rect 67222 481118 67306 481354
rect 67542 481118 102986 481354
rect 103222 481118 103306 481354
rect 103542 481118 138986 481354
rect 139222 481118 139306 481354
rect 139542 481118 174986 481354
rect 175222 481118 175306 481354
rect 175542 481118 210986 481354
rect 211222 481118 211306 481354
rect 211542 481118 246986 481354
rect 247222 481118 247306 481354
rect 247542 481118 282986 481354
rect 283222 481118 283306 481354
rect 283542 481118 283574 481354
rect 66954 481086 283574 481118
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect 63234 477954 279854 477986
rect 63234 477718 63266 477954
rect 63502 477718 63586 477954
rect 63822 477718 99266 477954
rect 99502 477718 99586 477954
rect 99822 477718 135266 477954
rect 135502 477718 135586 477954
rect 135822 477718 171266 477954
rect 171502 477718 171586 477954
rect 171822 477718 207266 477954
rect 207502 477718 207586 477954
rect 207822 477718 243266 477954
rect 243502 477718 243586 477954
rect 243822 477718 279266 477954
rect 279502 477718 279586 477954
rect 279822 477718 279854 477954
rect 63234 477634 279854 477718
rect 63234 477398 63266 477634
rect 63502 477398 63586 477634
rect 63822 477398 99266 477634
rect 99502 477398 99586 477634
rect 99822 477398 135266 477634
rect 135502 477398 135586 477634
rect 135822 477398 171266 477634
rect 171502 477398 171586 477634
rect 171822 477398 207266 477634
rect 207502 477398 207586 477634
rect 207822 477398 243266 477634
rect 243502 477398 243586 477634
rect 243822 477398 279266 477634
rect 279502 477398 279586 477634
rect 279822 477398 279854 477634
rect 63234 477366 279854 477398
rect 59514 476114 276134 476146
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 59514 475794 276134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 59514 475526 276134 475558
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect 91794 472394 272414 472426
rect 91794 472158 91826 472394
rect 92062 472158 92146 472394
rect 92382 472158 127826 472394
rect 128062 472158 128146 472394
rect 128382 472158 163826 472394
rect 164062 472158 164146 472394
rect 164382 472158 199826 472394
rect 200062 472158 200146 472394
rect 200382 472158 235826 472394
rect 236062 472158 236146 472394
rect 236382 472158 271826 472394
rect 272062 472158 272146 472394
rect 272382 472158 272414 472394
rect 91794 472074 272414 472158
rect 91794 471838 91826 472074
rect 92062 471838 92146 472074
rect 92382 471838 127826 472074
rect 128062 471838 128146 472074
rect 128382 471838 163826 472074
rect 164062 471838 164146 472074
rect 164382 471838 199826 472074
rect 200062 471838 200146 472074
rect 200382 471838 235826 472074
rect 236062 471838 236146 472074
rect 236382 471838 271826 472074
rect 272062 471838 272146 472074
rect 272382 471838 272414 472074
rect 91794 471806 272414 471838
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 380328 453454
rect 380564 453218 516056 453454
rect 516292 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 380328 453134
rect 380564 452898 516056 453134
rect 516292 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 381008 435454
rect 381244 435218 515376 435454
rect 515612 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 381008 435134
rect 381244 434898 515376 435134
rect 515612 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 380328 417454
rect 380564 417218 516056 417454
rect 516292 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 380328 417134
rect 380564 416898 516056 417134
rect 516292 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 61008 399454
rect 61244 399218 195376 399454
rect 195612 399218 221008 399454
rect 221244 399218 355376 399454
rect 355612 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 381008 399454
rect 381244 399218 515376 399454
rect 515612 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 61008 399134
rect 61244 398898 195376 399134
rect 195612 398898 221008 399134
rect 221244 398898 355376 399134
rect 355612 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 381008 399134
rect 381244 398898 515376 399134
rect 515612 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect 66954 373674 499574 373706
rect 66954 373438 66986 373674
rect 67222 373438 67306 373674
rect 67542 373438 102986 373674
rect 103222 373438 103306 373674
rect 103542 373438 138986 373674
rect 139222 373438 139306 373674
rect 139542 373438 174986 373674
rect 175222 373438 175306 373674
rect 175542 373438 210986 373674
rect 211222 373438 211306 373674
rect 211542 373438 246986 373674
rect 247222 373438 247306 373674
rect 247542 373438 282986 373674
rect 283222 373438 283306 373674
rect 283542 373438 318986 373674
rect 319222 373438 319306 373674
rect 319542 373438 354986 373674
rect 355222 373438 355306 373674
rect 355542 373438 390986 373674
rect 391222 373438 391306 373674
rect 391542 373438 426986 373674
rect 427222 373438 427306 373674
rect 427542 373438 462986 373674
rect 463222 373438 463306 373674
rect 463542 373438 498986 373674
rect 499222 373438 499306 373674
rect 499542 373438 499574 373674
rect 66954 373354 499574 373438
rect 66954 373118 66986 373354
rect 67222 373118 67306 373354
rect 67542 373118 102986 373354
rect 103222 373118 103306 373354
rect 103542 373118 138986 373354
rect 139222 373118 139306 373354
rect 139542 373118 174986 373354
rect 175222 373118 175306 373354
rect 175542 373118 210986 373354
rect 211222 373118 211306 373354
rect 211542 373118 246986 373354
rect 247222 373118 247306 373354
rect 247542 373118 282986 373354
rect 283222 373118 283306 373354
rect 283542 373118 318986 373354
rect 319222 373118 319306 373354
rect 319542 373118 354986 373354
rect 355222 373118 355306 373354
rect 355542 373118 390986 373354
rect 391222 373118 391306 373354
rect 391542 373118 426986 373354
rect 427222 373118 427306 373354
rect 427542 373118 462986 373354
rect 463222 373118 463306 373354
rect 463542 373118 498986 373354
rect 499222 373118 499306 373354
rect 499542 373118 499574 373354
rect 66954 373086 499574 373118
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect 63234 369954 495854 369986
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 63234 369634 495854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 63234 369366 495854 369398
rect 59514 368114 492134 368146
rect 59514 367878 59546 368114
rect 59782 367878 59866 368114
rect 60102 367878 95546 368114
rect 95782 367878 95866 368114
rect 96102 367878 131546 368114
rect 131782 367878 131866 368114
rect 132102 367878 167546 368114
rect 167782 367878 167866 368114
rect 168102 367878 203546 368114
rect 203782 367878 203866 368114
rect 204102 367878 239546 368114
rect 239782 367878 239866 368114
rect 240102 367878 275546 368114
rect 275782 367878 275866 368114
rect 276102 367878 311546 368114
rect 311782 367878 311866 368114
rect 312102 367878 347546 368114
rect 347782 367878 347866 368114
rect 348102 367878 383546 368114
rect 383782 367878 383866 368114
rect 384102 367878 419546 368114
rect 419782 367878 419866 368114
rect 420102 367878 455546 368114
rect 455782 367878 455866 368114
rect 456102 367878 491546 368114
rect 491782 367878 491866 368114
rect 492102 367878 492134 368114
rect 59514 367794 492134 367878
rect 59514 367558 59546 367794
rect 59782 367558 59866 367794
rect 60102 367558 95546 367794
rect 95782 367558 95866 367794
rect 96102 367558 131546 367794
rect 131782 367558 131866 367794
rect 132102 367558 167546 367794
rect 167782 367558 167866 367794
rect 168102 367558 203546 367794
rect 203782 367558 203866 367794
rect 204102 367558 239546 367794
rect 239782 367558 239866 367794
rect 240102 367558 275546 367794
rect 275782 367558 275866 367794
rect 276102 367558 311546 367794
rect 311782 367558 311866 367794
rect 312102 367558 347546 367794
rect 347782 367558 347866 367794
rect 348102 367558 383546 367794
rect 383782 367558 383866 367794
rect 384102 367558 419546 367794
rect 419782 367558 419866 367794
rect 420102 367558 455546 367794
rect 455782 367558 455866 367794
rect 456102 367558 491546 367794
rect 491782 367558 491866 367794
rect 492102 367558 492134 367794
rect 59514 367526 492134 367558
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect 91794 364394 488414 364426
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 91794 364074 488414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 91794 363806 488414 363838
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 60328 345454
rect 60564 345218 196056 345454
rect 196292 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 220328 345454
rect 220564 345218 356056 345454
rect 356292 345218 380328 345454
rect 380564 345218 516056 345454
rect 516292 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 60328 345134
rect 60564 344898 196056 345134
rect 196292 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 220328 345134
rect 220564 344898 356056 345134
rect 356292 344898 380328 345134
rect 380564 344898 516056 345134
rect 516292 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 61008 327454
rect 61244 327218 195376 327454
rect 195612 327218 221008 327454
rect 221244 327218 355376 327454
rect 355612 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 381008 327454
rect 381244 327218 515376 327454
rect 515612 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 61008 327134
rect 61244 326898 195376 327134
rect 195612 326898 221008 327134
rect 221244 326898 355376 327134
rect 355612 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 381008 327134
rect 381244 326898 515376 327134
rect 515612 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 60328 309454
rect 60564 309218 196056 309454
rect 196292 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 220328 309454
rect 220564 309218 356056 309454
rect 356292 309218 380328 309454
rect 380564 309218 516056 309454
rect 516292 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 60328 309134
rect 60564 308898 196056 309134
rect 196292 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 220328 309134
rect 220564 308898 356056 309134
rect 356292 308898 380328 309134
rect 380564 308898 516056 309134
rect 516292 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 61008 291454
rect 61244 291218 195376 291454
rect 195612 291218 221008 291454
rect 221244 291218 355376 291454
rect 355612 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 381008 291454
rect 381244 291218 515376 291454
rect 515612 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 61008 291134
rect 61244 290898 195376 291134
rect 195612 290898 221008 291134
rect 221244 290898 355376 291134
rect 355612 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 381008 291134
rect 381244 290898 515376 291134
rect 515612 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect 66954 265674 499574 265706
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 66954 265354 499574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 66954 265086 499574 265118
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect 63234 261954 495854 261986
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 63234 261634 495854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 63234 261366 495854 261398
rect 59514 260114 492134 260146
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 59514 259794 492134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 59514 259526 492134 259558
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect 91794 256394 488414 256426
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 91794 256074 488414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 91794 255806 488414 255838
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 60328 237454
rect 60564 237218 196056 237454
rect 196292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 220328 237454
rect 220564 237218 356056 237454
rect 356292 237218 380328 237454
rect 380564 237218 516056 237454
rect 516292 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 60328 237134
rect 60564 236898 196056 237134
rect 196292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 220328 237134
rect 220564 236898 356056 237134
rect 356292 236898 380328 237134
rect 380564 236898 516056 237134
rect 516292 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 61008 219454
rect 61244 219218 195376 219454
rect 195612 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 381008 219454
rect 381244 219218 515376 219454
rect 515612 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 61008 219134
rect 61244 218898 195376 219134
rect 195612 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 381008 219134
rect 381244 218898 515376 219134
rect 515612 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 60328 201454
rect 60564 201218 196056 201454
rect 196292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 220328 201454
rect 220564 201218 356056 201454
rect 356292 201218 380328 201454
rect 380564 201218 516056 201454
rect 516292 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 60328 201134
rect 60564 200898 196056 201134
rect 196292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 220328 201134
rect 220564 200898 356056 201134
rect 356292 200898 380328 201134
rect 380564 200898 516056 201134
rect 516292 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 61008 183454
rect 61244 183218 195376 183454
rect 195612 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 381008 183454
rect 381244 183218 515376 183454
rect 515612 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 61008 183134
rect 61244 182898 195376 183134
rect 195612 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 381008 183134
rect 381244 182898 515376 183134
rect 515612 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect 66954 157674 499574 157706
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 66954 157354 499574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 66954 157086 499574 157118
rect 63234 155834 495854 155866
rect 63234 155598 63266 155834
rect 63502 155598 63586 155834
rect 63822 155598 99266 155834
rect 99502 155598 99586 155834
rect 99822 155598 135266 155834
rect 135502 155598 135586 155834
rect 135822 155598 171266 155834
rect 171502 155598 171586 155834
rect 171822 155598 207266 155834
rect 207502 155598 207586 155834
rect 207822 155598 243266 155834
rect 243502 155598 243586 155834
rect 243822 155598 279266 155834
rect 279502 155598 279586 155834
rect 279822 155598 315266 155834
rect 315502 155598 315586 155834
rect 315822 155598 351266 155834
rect 351502 155598 351586 155834
rect 351822 155598 387266 155834
rect 387502 155598 387586 155834
rect 387822 155598 423266 155834
rect 423502 155598 423586 155834
rect 423822 155598 459266 155834
rect 459502 155598 459586 155834
rect 459822 155598 495266 155834
rect 495502 155598 495586 155834
rect 495822 155598 495854 155834
rect 63234 155514 495854 155598
rect 63234 155278 63266 155514
rect 63502 155278 63586 155514
rect 63822 155278 99266 155514
rect 99502 155278 99586 155514
rect 99822 155278 135266 155514
rect 135502 155278 135586 155514
rect 135822 155278 171266 155514
rect 171502 155278 171586 155514
rect 171822 155278 207266 155514
rect 207502 155278 207586 155514
rect 207822 155278 243266 155514
rect 243502 155278 243586 155514
rect 243822 155278 279266 155514
rect 279502 155278 279586 155514
rect 279822 155278 315266 155514
rect 315502 155278 315586 155514
rect 315822 155278 351266 155514
rect 351502 155278 351586 155514
rect 351822 155278 387266 155514
rect 387502 155278 387586 155514
rect 387822 155278 423266 155514
rect 423502 155278 423586 155514
rect 423822 155278 459266 155514
rect 459502 155278 459586 155514
rect 459822 155278 495266 155514
rect 495502 155278 495586 155514
rect 495822 155278 495854 155514
rect 63234 155246 495854 155278
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect 59514 152114 492134 152146
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 59514 151794 492134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 59514 151526 492134 151558
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect 91794 148394 488414 148426
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 91794 148074 488414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 91794 147806 488414 147838
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 60328 129454
rect 60564 129218 196056 129454
rect 196292 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 220328 129454
rect 220564 129218 356056 129454
rect 356292 129218 380328 129454
rect 380564 129218 516056 129454
rect 516292 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 60328 129134
rect 60564 128898 196056 129134
rect 196292 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 220328 129134
rect 220564 128898 356056 129134
rect 356292 128898 380328 129134
rect 380564 128898 516056 129134
rect 516292 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 61008 111454
rect 61244 111218 195376 111454
rect 195612 111218 221008 111454
rect 221244 111218 355376 111454
rect 355612 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 381008 111454
rect 381244 111218 515376 111454
rect 515612 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 61008 111134
rect 61244 110898 195376 111134
rect 195612 110898 221008 111134
rect 221244 110898 355376 111134
rect 355612 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 381008 111134
rect 381244 110898 515376 111134
rect 515612 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 60328 93454
rect 60564 93218 196056 93454
rect 196292 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 220328 93454
rect 220564 93218 356056 93454
rect 356292 93218 380328 93454
rect 380564 93218 516056 93454
rect 516292 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 60328 93134
rect 60564 92898 196056 93134
rect 196292 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 220328 93134
rect 220564 92898 356056 93134
rect 356292 92898 380328 93134
rect 380564 92898 516056 93134
rect 516292 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 61008 75454
rect 61244 75218 195376 75454
rect 195612 75218 221008 75454
rect 221244 75218 355376 75454
rect 355612 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 381008 75454
rect 381244 75218 515376 75454
rect 515612 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 61008 75134
rect 61244 74898 195376 75134
rect 195612 74898 221008 75134
rect 221244 74898 355376 75134
rect 355612 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 381008 75134
rect 381244 74898 515376 75134
rect 515612 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst1
timestamp 0
transform 1 0 60000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst2
timestamp 0
transform 1 0 60000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst0
timestamp 0
transform 1 0 380000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst1
timestamp 0
transform 1 0 380000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst2
timestamp 0
transform 1 0 380000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst3
timestamp 0
transform 1 0 380000 0 1 381000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 381000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst1
timestamp 0
transform 1 0 220000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst2
timestamp 0
transform 1 0 220000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst3
timestamp 0
transform 1 0 220000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst4
timestamp 0
transform 1 0 220000 0 1 381000
box 0 0 136620 83308
use VerySimpleCPU_core  inst_agent_1
timestamp 0
transform 1 0 60000 0 1 568000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_codemaker
timestamp 0
transform 1 0 240000 0 1 568000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_control_tower
timestamp 0
transform 1 0 150000 0 1 568000
box 0 0 60955 63099
use main_controller  inst_main_controller
timestamp 0
transform 1 0 60000 0 1 488000
box 0 0 240000 60000
use main_memory  inst_main_memory
timestamp 0
transform 1 0 325000 0 1 522000
box 0 0 108889 111033
use uart  inst_uart
timestamp 0
transform 1 0 460000 0 1 578000
box 0 0 50000 50000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s 73794 559926 290414 560546 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 145308 74414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 145308 110414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 145308 146414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 145308 182414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 145308 218414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 145308 254414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 145308 290414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 145308 326414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 145308 398414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 145308 434414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 145308 470414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 145308 506414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 252308 74414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 252308 110414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 252308 146414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 252308 182414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 252308 218414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 252308 254414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 252308 290414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 252308 326414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 252308 398414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 252308 434414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 252308 470414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 252308 506414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 359308 74414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 359308 110414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 359308 146414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 359308 182414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 359308 218414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 359308 254414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 359308 290414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 359308 326414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 359308 398414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 359308 434414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 359308 470414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 359308 506414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 466308 74414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 466308 110414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 466308 146414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 466308 182414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 466308 218414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 466308 254414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 466308 290414 486000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 466308 326414 520000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 520000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 466308 398414 520000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 466308 434414 520000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 550000 74414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 550000 110414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 550000 182414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 550000 254414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 550000 290414 566000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 466308 470414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 466308 506414 576000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 633099 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 633099 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 550000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 633099 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 550000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 633099 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 633099 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 635033 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 635033 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 635033 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 635033 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 630000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 630000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s 77514 563646 294134 564266 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 145308 78134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 145308 114134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 145308 150134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 145308 186134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 145308 222134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 145308 258134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 145308 294134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 145308 330134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 145308 402134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 145308 438134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 145308 474134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 145308 510134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 252308 78134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 252308 114134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 252308 150134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 252308 186134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 252308 222134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 252308 258134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 252308 294134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 252308 330134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 252308 402134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 252308 438134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 252308 474134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 252308 510134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 359308 78134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 359308 114134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 359308 150134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 359308 186134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 359308 222134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 359308 258134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 359308 294134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 359308 330134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 359308 402134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 359308 438134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 359308 474134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 359308 510134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 466308 78134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 466308 114134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 466308 150134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 466308 186134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 466308 222134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 466308 258134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 466308 294134 486000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 466308 330134 520000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 520000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 466308 402134 520000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 550000 78134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 550000 114134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 550000 150134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 550000 186134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 550000 258134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 550000 294134 566000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 466308 474134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 466308 510134 576000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 633099 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 633099 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 633099 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 633099 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 550000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 633099 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 633099 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 635033 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 635033 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 635033 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 466308 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 630000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 630000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 145308 81854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 145308 117854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 145308 153854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 145308 189854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 145308 225854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 145308 261854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 145308 297854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 145308 333854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 145308 405854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 145308 441854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 145308 477854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 145308 513854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 252308 81854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 252308 117854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 252308 153854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 252308 189854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 252308 225854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 252308 261854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 252308 297854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 252308 333854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 252308 405854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 252308 441854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 252308 477854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 252308 513854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 359308 81854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 359308 117854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 359308 153854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 359308 189854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 359308 225854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 359308 261854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 359308 297854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 359308 333854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 359308 405854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 359308 441854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 359308 477854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 359308 513854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 466308 81854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 466308 117854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 466308 153854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 466308 189854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 466308 225854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 466308 261854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 466308 297854 486000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 466308 333854 520000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 520000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 466308 405854 520000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 550000 81854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 550000 117854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 550000 153854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 550000 189854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 550000 261854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 550000 297854 566000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 466308 477854 576000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 633099 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 633099 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 633099 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 633099 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 550000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 633099 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 633099 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 635033 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 635033 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 635033 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 466308 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 630000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 466308 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 145308 85574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 145308 121574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 145308 157574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 145308 193574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 145308 229574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 145308 265574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 145308 301574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 145308 337574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 145308 409574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 145308 445574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 145308 481574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 145308 517574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 252308 85574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 252308 121574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 252308 157574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 252308 193574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 252308 229574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 252308 265574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 252308 301574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 252308 337574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 252308 409574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 252308 445574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 252308 481574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 252308 517574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 359308 85574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 359308 121574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 359308 157574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 359308 193574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 359308 229574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 359308 265574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 359308 301574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 359308 337574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 359308 409574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 359308 445574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 359308 481574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 359308 517574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 466308 85574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 466308 121574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 466308 157574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 466308 193574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 466308 229574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 466308 265574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 466308 301574 486000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 466308 337574 520000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 520000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 466308 409574 520000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 550000 85574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 550000 121574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 550000 157574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 550000 193574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 550000 265574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 550000 301574 566000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 466308 481574 576000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 633099 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 633099 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 633099 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 633099 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 550000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 633099 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 633099 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 635033 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 635033 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 635033 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 466308 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 630000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 466308 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 155246 495854 155866 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 261366 495854 261986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 369366 495854 369986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 477366 279854 477986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 551246 279854 551866 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 145308 63854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 145308 99854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 145308 135854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 145308 171854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 145308 243854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 145308 279854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 145308 315854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 145308 351854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 145308 387854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 145308 423854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 145308 459854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 145308 495854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 252308 63854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 252308 99854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 252308 135854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 252308 171854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 252308 243854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 252308 279854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 252308 315854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 252308 351854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 252308 387854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 252308 423854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 252308 459854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 252308 495854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 359308 63854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 359308 99854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 359308 135854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 359308 171854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 359308 243854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 359308 279854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 359308 315854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 359308 351854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 359308 387854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 359308 423854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 359308 459854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 359308 495854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 466308 63854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 466308 99854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 466308 135854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 466308 171854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 466308 243854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 466308 279854 486000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 466308 351854 520000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 466308 387854 520000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 466308 423854 520000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 550000 63854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 550000 99854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 550000 171854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 550000 207854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 550000 243854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 550000 279854 566000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 466308 459854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 466308 495854 576000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 633099 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 633099 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 550000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 633099 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 633099 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 633099 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 633099 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 466308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 635033 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 635033 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 635033 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 630000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 630000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 157086 499574 157706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 265086 499574 265706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 373086 499574 373706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 481086 283574 481706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 554966 283574 555586 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 145308 67574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 145308 103574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 145308 139574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 145308 175574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 145308 247574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 145308 283574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 145308 319574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 145308 355574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 145308 391574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 145308 427574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 145308 463574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 145308 499574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 252308 67574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 252308 103574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 252308 139574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 252308 175574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 252308 247574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 252308 283574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 252308 319574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 252308 355574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 252308 391574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 252308 427574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 252308 463574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 252308 499574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 359308 67574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 359308 103574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 359308 139574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 359308 175574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 359308 247574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 359308 283574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 359308 319574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 359308 355574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 359308 391574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 359308 427574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 359308 463574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 359308 499574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 466308 67574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 466308 103574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 466308 139574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 466308 175574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 466308 247574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 466308 283574 486000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 466308 355574 520000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 466308 391574 520000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 466308 427574 520000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 550000 67574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 550000 103574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 550000 175574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 550000 211574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 550000 247574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 550000 283574 566000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 466308 463574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 466308 499574 576000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 633099 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 633099 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 550000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 633099 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 633099 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 633099 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 633099 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 466308 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 635033 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 635033 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 635033 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 630000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 630000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 147806 488414 148426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 255806 488414 256426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 363806 488414 364426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 471806 272414 472426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 145308 92414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 145308 128414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 145308 164414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 145308 236414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 145308 272414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 145308 308414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 145308 344414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 145308 380414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 145308 416414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 145308 452414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 145308 488414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 252308 92414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 252308 128414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 252308 164414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 252308 236414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 252308 272414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 252308 308414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 252308 344414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 252308 380414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 252308 416414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 252308 452414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 252308 488414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 359308 92414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 359308 128414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 359308 164414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 359308 236414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 359308 272414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 359308 308414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 359308 344414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 359308 380414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 359308 416414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 359308 452414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 359308 488414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 466308 92414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 466308 128414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 466308 164414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 466308 236414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 466308 272414 486000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 466308 344414 520000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 466308 380414 520000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 466308 416414 520000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 550000 92414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 550000 164414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 550000 200414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 550000 272414 566000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 466308 488414 576000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 633099 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 550000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 633099 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 633099 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 550000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 633099 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 466308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 635033 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 635033 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 635033 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 466308 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 630000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 151526 492134 152146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 259526 492134 260146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 367526 492134 368146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 475526 276134 476146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 145308 60134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 145308 96134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 145308 132134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 145308 168134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 145308 240134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 145308 276134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 145308 312134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 145308 348134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 145308 384134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 145308 420134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 145308 456134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 145308 492134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 252308 60134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 252308 96134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 252308 132134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 252308 168134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 252308 240134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 252308 276134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 252308 312134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 252308 348134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 252308 384134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 252308 420134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 252308 456134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 252308 492134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 359308 60134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 359308 96134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 359308 132134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 359308 168134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 359308 240134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 359308 276134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 359308 312134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 359308 348134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 359308 384134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 359308 420134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 359308 456134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 359308 492134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 466308 60134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 466308 96134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 466308 132134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 466308 168134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 466308 240134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 466308 276134 486000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 466308 348134 520000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 466308 384134 520000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 466308 420134 520000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 550000 60134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 550000 96134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 550000 168134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 550000 204134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 550000 240134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 550000 276134 566000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 466308 492134 576000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 633099 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 633099 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 550000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 633099 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 633099 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 633099 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 633099 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 466308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 635033 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 635033 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 635033 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 466308 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 630000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
