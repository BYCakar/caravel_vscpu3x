VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO uart
  CLASS BLOCK ;
  FOREIGN uart ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END clk
  PIN dvsr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 246.000 235.430 250.000 ;
    END
  END dvsr[0]
  PIN dvsr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END dvsr[1]
  PIN dvsr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 246.000 87.310 250.000 ;
    END
  END dvsr[2]
  PIN dvsr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END dvsr[3]
  PIN dvsr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 78.240 250.000 78.840 ;
    END
  END dvsr[4]
  PIN dvsr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 246.000 145.270 250.000 ;
    END
  END dvsr[5]
  PIN dvsr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END dvsr[6]
  PIN dvsr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 139.440 250.000 140.040 ;
    END
  END dvsr[7]
  PIN r_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END r_data[0]
  PIN r_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 170.040 250.000 170.640 ;
    END
  END r_data[1]
  PIN r_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END r_data[2]
  PIN r_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END r_data[3]
  PIN r_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 246.000 174.250 250.000 ;
    END
  END r_data[4]
  PIN r_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 246.000 206.450 250.000 ;
    END
  END r_data[5]
  PIN r_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END r_data[6]
  PIN r_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 246.000 58.330 250.000 ;
    END
  END r_data[7]
  PIN rd_uart
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END rd_uart
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END reset
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 13.640 250.000 14.240 ;
    END
  END rx
  PIN rx_empty
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END rx_empty
  PIN rx_fifo_flush_enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END rx_fifo_flush_enable
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 246.000 26.130 250.000 ;
    END
  END tx
  PIN tx_full
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 47.640 250.000 48.240 ;
    END
  END tx_full
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
  END vssd1
  PIN w_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END w_data[0]
  PIN w_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 204.040 250.000 204.640 ;
    END
  END w_data[1]
  PIN w_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 234.640 250.000 235.240 ;
    END
  END w_data[2]
  PIN w_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END w_data[3]
  PIN w_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 246.000 116.290 250.000 ;
    END
  END w_data[4]
  PIN w_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END w_data[5]
  PIN w_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END w_data[6]
  PIN w_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END w_data[7]
  PIN wr_uart
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 246.000 108.840 250.000 109.440 ;
    END
  END wr_uart
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 0.070 10.240 244.260 236.880 ;
      LAYER met2 ;
        RECT 0.100 245.720 25.570 248.725 ;
        RECT 26.410 245.720 57.770 248.725 ;
        RECT 58.610 245.720 86.750 248.725 ;
        RECT 87.590 245.720 115.730 248.725 ;
        RECT 116.570 245.720 144.710 248.725 ;
        RECT 145.550 245.720 173.690 248.725 ;
        RECT 174.530 245.720 205.890 248.725 ;
        RECT 206.730 245.720 234.870 248.725 ;
        RECT 235.710 245.720 240.490 248.725 ;
        RECT 0.100 4.280 240.490 245.720 ;
        RECT 0.650 4.000 28.790 4.280 ;
        RECT 29.630 4.000 57.770 4.280 ;
        RECT 58.610 4.000 86.750 4.280 ;
        RECT 87.590 4.000 115.730 4.280 ;
        RECT 116.570 4.000 147.930 4.280 ;
        RECT 148.770 4.000 176.910 4.280 ;
        RECT 177.750 4.000 205.890 4.280 ;
        RECT 206.730 4.000 234.870 4.280 ;
        RECT 235.710 4.000 240.490 4.280 ;
      LAYER met3 ;
        RECT 4.400 247.840 246.000 248.705 ;
        RECT 4.000 235.640 246.000 247.840 ;
        RECT 4.000 234.240 245.600 235.640 ;
        RECT 4.000 218.640 246.000 234.240 ;
        RECT 4.400 217.240 246.000 218.640 ;
        RECT 4.000 205.040 246.000 217.240 ;
        RECT 4.000 203.640 245.600 205.040 ;
        RECT 4.000 188.040 246.000 203.640 ;
        RECT 4.400 186.640 246.000 188.040 ;
        RECT 4.000 171.040 246.000 186.640 ;
        RECT 4.000 169.640 245.600 171.040 ;
        RECT 4.000 157.440 246.000 169.640 ;
        RECT 4.400 156.040 246.000 157.440 ;
        RECT 4.000 140.440 246.000 156.040 ;
        RECT 4.000 139.040 245.600 140.440 ;
        RECT 4.000 123.440 246.000 139.040 ;
        RECT 4.400 122.040 246.000 123.440 ;
        RECT 4.000 109.840 246.000 122.040 ;
        RECT 4.000 108.440 245.600 109.840 ;
        RECT 4.000 92.840 246.000 108.440 ;
        RECT 4.400 91.440 246.000 92.840 ;
        RECT 4.000 79.240 246.000 91.440 ;
        RECT 4.000 77.840 245.600 79.240 ;
        RECT 4.000 62.240 246.000 77.840 ;
        RECT 4.400 60.840 246.000 62.240 ;
        RECT 4.000 48.640 246.000 60.840 ;
        RECT 4.000 47.240 245.600 48.640 ;
        RECT 4.000 31.640 246.000 47.240 ;
        RECT 4.400 30.240 246.000 31.640 ;
        RECT 4.000 14.640 246.000 30.240 ;
        RECT 4.000 13.240 245.600 14.640 ;
        RECT 4.000 10.715 246.000 13.240 ;
  END
END uart
END LIBRARY

